magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 3442 582
<< pwell >>
rect 1 177 185 203
rect 735 177 1013 203
rect 1563 177 1841 203
rect 2391 177 2669 203
rect 3219 177 3403 203
rect 1 21 3403 177
rect 29 -17 63 21
rect 857 -17 891 21
rect 1685 -17 1719 21
rect 2513 -17 2547 21
rect 3341 -17 3375 21
<< scnmos >>
rect 79 47 109 177
rect 174 47 204 151
rect 387 47 417 151
rect 503 47 533 151
rect 716 47 746 151
rect 811 47 841 177
rect 907 47 937 177
rect 1002 47 1032 151
rect 1215 47 1245 151
rect 1331 47 1361 151
rect 1544 47 1574 151
rect 1639 47 1669 177
rect 1735 47 1765 177
rect 1830 47 1860 151
rect 2043 47 2073 151
rect 2159 47 2189 151
rect 2372 47 2402 151
rect 2467 47 2497 177
rect 2563 47 2593 177
rect 2658 47 2688 151
rect 2871 47 2901 151
rect 2987 47 3017 151
rect 3200 47 3230 151
rect 3295 47 3325 177
<< scpmoshvt >>
rect 81 297 117 497
rect 186 333 222 497
rect 384 297 420 497
rect 500 297 536 497
rect 698 333 734 497
rect 803 297 839 497
rect 909 297 945 497
rect 1014 333 1050 497
rect 1212 297 1248 497
rect 1328 297 1364 497
rect 1526 333 1562 497
rect 1631 297 1667 497
rect 1737 297 1773 497
rect 1842 333 1878 497
rect 2040 297 2076 497
rect 2156 297 2192 497
rect 2354 333 2390 497
rect 2459 297 2495 497
rect 2565 297 2601 497
rect 2670 333 2706 497
rect 2868 297 2904 497
rect 2984 297 3020 497
rect 3182 333 3218 497
rect 3287 297 3323 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 151 159 177
rect 761 151 811 177
rect 109 47 174 151
rect 204 116 256 151
rect 204 82 214 116
rect 248 82 256 116
rect 204 47 256 82
rect 330 116 387 151
rect 330 82 338 116
rect 372 82 387 116
rect 330 47 387 82
rect 417 116 503 151
rect 417 82 443 116
rect 477 82 503 116
rect 417 47 503 82
rect 533 116 590 151
rect 533 82 548 116
rect 582 82 590 116
rect 533 47 590 82
rect 664 116 716 151
rect 664 82 672 116
rect 706 82 716 116
rect 664 47 716 82
rect 746 47 811 151
rect 841 161 907 177
rect 841 127 857 161
rect 891 127 907 161
rect 841 93 907 127
rect 841 59 857 93
rect 891 59 907 93
rect 841 47 907 59
rect 937 151 987 177
rect 1589 151 1639 177
rect 937 47 1002 151
rect 1032 116 1084 151
rect 1032 82 1042 116
rect 1076 82 1084 116
rect 1032 47 1084 82
rect 1158 116 1215 151
rect 1158 82 1166 116
rect 1200 82 1215 116
rect 1158 47 1215 82
rect 1245 116 1331 151
rect 1245 82 1271 116
rect 1305 82 1331 116
rect 1245 47 1331 82
rect 1361 116 1418 151
rect 1361 82 1376 116
rect 1410 82 1418 116
rect 1361 47 1418 82
rect 1492 116 1544 151
rect 1492 82 1500 116
rect 1534 82 1544 116
rect 1492 47 1544 82
rect 1574 47 1639 151
rect 1669 161 1735 177
rect 1669 127 1685 161
rect 1719 127 1735 161
rect 1669 93 1735 127
rect 1669 59 1685 93
rect 1719 59 1735 93
rect 1669 47 1735 59
rect 1765 151 1815 177
rect 2417 151 2467 177
rect 1765 47 1830 151
rect 1860 116 1912 151
rect 1860 82 1870 116
rect 1904 82 1912 116
rect 1860 47 1912 82
rect 1986 116 2043 151
rect 1986 82 1994 116
rect 2028 82 2043 116
rect 1986 47 2043 82
rect 2073 116 2159 151
rect 2073 82 2099 116
rect 2133 82 2159 116
rect 2073 47 2159 82
rect 2189 116 2246 151
rect 2189 82 2204 116
rect 2238 82 2246 116
rect 2189 47 2246 82
rect 2320 116 2372 151
rect 2320 82 2328 116
rect 2362 82 2372 116
rect 2320 47 2372 82
rect 2402 47 2467 151
rect 2497 161 2563 177
rect 2497 127 2513 161
rect 2547 127 2563 161
rect 2497 93 2563 127
rect 2497 59 2513 93
rect 2547 59 2563 93
rect 2497 47 2563 59
rect 2593 151 2643 177
rect 3245 151 3295 177
rect 2593 47 2658 151
rect 2688 116 2740 151
rect 2688 82 2698 116
rect 2732 82 2740 116
rect 2688 47 2740 82
rect 2814 116 2871 151
rect 2814 82 2822 116
rect 2856 82 2871 116
rect 2814 47 2871 82
rect 2901 116 2987 151
rect 2901 82 2927 116
rect 2961 82 2987 116
rect 2901 47 2987 82
rect 3017 116 3074 151
rect 3017 82 3032 116
rect 3066 82 3074 116
rect 3017 47 3074 82
rect 3148 116 3200 151
rect 3148 82 3156 116
rect 3190 82 3200 116
rect 3148 47 3200 82
rect 3230 47 3295 151
rect 3325 161 3377 177
rect 3325 127 3335 161
rect 3369 127 3377 161
rect 3325 93 3377 127
rect 3325 59 3335 93
rect 3369 59 3377 93
rect 3325 47 3377 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 333 186 497
rect 222 485 276 497
rect 222 451 234 485
rect 268 451 276 485
rect 222 417 276 451
rect 222 383 234 417
rect 268 383 276 417
rect 222 333 276 383
rect 330 479 384 497
rect 330 445 338 479
rect 372 445 384 479
rect 330 411 384 445
rect 330 377 338 411
rect 372 377 384 411
rect 330 343 384 377
rect 117 297 169 333
rect 330 309 338 343
rect 372 309 384 343
rect 330 297 384 309
rect 420 479 500 497
rect 420 445 443 479
rect 477 445 500 479
rect 420 411 500 445
rect 420 377 443 411
rect 477 377 500 411
rect 420 343 500 377
rect 420 309 443 343
rect 477 309 500 343
rect 420 297 500 309
rect 536 479 590 497
rect 536 445 548 479
rect 582 445 590 479
rect 536 411 590 445
rect 536 377 548 411
rect 582 377 590 411
rect 536 343 590 377
rect 536 309 548 343
rect 582 309 590 343
rect 644 485 698 497
rect 644 451 652 485
rect 686 451 698 485
rect 644 417 698 451
rect 644 383 652 417
rect 686 383 698 417
rect 644 333 698 383
rect 734 333 803 497
rect 536 297 590 309
rect 751 297 803 333
rect 839 485 909 497
rect 839 451 857 485
rect 891 451 909 485
rect 839 417 909 451
rect 839 383 857 417
rect 891 383 909 417
rect 839 349 909 383
rect 839 315 857 349
rect 891 315 909 349
rect 839 297 909 315
rect 945 333 1014 497
rect 1050 485 1104 497
rect 1050 451 1062 485
rect 1096 451 1104 485
rect 1050 417 1104 451
rect 1050 383 1062 417
rect 1096 383 1104 417
rect 1050 333 1104 383
rect 1158 479 1212 497
rect 1158 445 1166 479
rect 1200 445 1212 479
rect 1158 411 1212 445
rect 1158 377 1166 411
rect 1200 377 1212 411
rect 1158 343 1212 377
rect 945 297 997 333
rect 1158 309 1166 343
rect 1200 309 1212 343
rect 1158 297 1212 309
rect 1248 479 1328 497
rect 1248 445 1271 479
rect 1305 445 1328 479
rect 1248 411 1328 445
rect 1248 377 1271 411
rect 1305 377 1328 411
rect 1248 343 1328 377
rect 1248 309 1271 343
rect 1305 309 1328 343
rect 1248 297 1328 309
rect 1364 479 1418 497
rect 1364 445 1376 479
rect 1410 445 1418 479
rect 1364 411 1418 445
rect 1364 377 1376 411
rect 1410 377 1418 411
rect 1364 343 1418 377
rect 1364 309 1376 343
rect 1410 309 1418 343
rect 1472 485 1526 497
rect 1472 451 1480 485
rect 1514 451 1526 485
rect 1472 417 1526 451
rect 1472 383 1480 417
rect 1514 383 1526 417
rect 1472 333 1526 383
rect 1562 333 1631 497
rect 1364 297 1418 309
rect 1579 297 1631 333
rect 1667 485 1737 497
rect 1667 451 1685 485
rect 1719 451 1737 485
rect 1667 417 1737 451
rect 1667 383 1685 417
rect 1719 383 1737 417
rect 1667 349 1737 383
rect 1667 315 1685 349
rect 1719 315 1737 349
rect 1667 297 1737 315
rect 1773 333 1842 497
rect 1878 485 1932 497
rect 1878 451 1890 485
rect 1924 451 1932 485
rect 1878 417 1932 451
rect 1878 383 1890 417
rect 1924 383 1932 417
rect 1878 333 1932 383
rect 1986 479 2040 497
rect 1986 445 1994 479
rect 2028 445 2040 479
rect 1986 411 2040 445
rect 1986 377 1994 411
rect 2028 377 2040 411
rect 1986 343 2040 377
rect 1773 297 1825 333
rect 1986 309 1994 343
rect 2028 309 2040 343
rect 1986 297 2040 309
rect 2076 479 2156 497
rect 2076 445 2099 479
rect 2133 445 2156 479
rect 2076 411 2156 445
rect 2076 377 2099 411
rect 2133 377 2156 411
rect 2076 343 2156 377
rect 2076 309 2099 343
rect 2133 309 2156 343
rect 2076 297 2156 309
rect 2192 479 2246 497
rect 2192 445 2204 479
rect 2238 445 2246 479
rect 2192 411 2246 445
rect 2192 377 2204 411
rect 2238 377 2246 411
rect 2192 343 2246 377
rect 2192 309 2204 343
rect 2238 309 2246 343
rect 2300 485 2354 497
rect 2300 451 2308 485
rect 2342 451 2354 485
rect 2300 417 2354 451
rect 2300 383 2308 417
rect 2342 383 2354 417
rect 2300 333 2354 383
rect 2390 333 2459 497
rect 2192 297 2246 309
rect 2407 297 2459 333
rect 2495 485 2565 497
rect 2495 451 2513 485
rect 2547 451 2565 485
rect 2495 417 2565 451
rect 2495 383 2513 417
rect 2547 383 2565 417
rect 2495 349 2565 383
rect 2495 315 2513 349
rect 2547 315 2565 349
rect 2495 297 2565 315
rect 2601 333 2670 497
rect 2706 485 2760 497
rect 2706 451 2718 485
rect 2752 451 2760 485
rect 2706 417 2760 451
rect 2706 383 2718 417
rect 2752 383 2760 417
rect 2706 333 2760 383
rect 2814 479 2868 497
rect 2814 445 2822 479
rect 2856 445 2868 479
rect 2814 411 2868 445
rect 2814 377 2822 411
rect 2856 377 2868 411
rect 2814 343 2868 377
rect 2601 297 2653 333
rect 2814 309 2822 343
rect 2856 309 2868 343
rect 2814 297 2868 309
rect 2904 479 2984 497
rect 2904 445 2927 479
rect 2961 445 2984 479
rect 2904 411 2984 445
rect 2904 377 2927 411
rect 2961 377 2984 411
rect 2904 343 2984 377
rect 2904 309 2927 343
rect 2961 309 2984 343
rect 2904 297 2984 309
rect 3020 479 3074 497
rect 3020 445 3032 479
rect 3066 445 3074 479
rect 3020 411 3074 445
rect 3020 377 3032 411
rect 3066 377 3074 411
rect 3020 343 3074 377
rect 3020 309 3032 343
rect 3066 309 3074 343
rect 3128 485 3182 497
rect 3128 451 3136 485
rect 3170 451 3182 485
rect 3128 417 3182 451
rect 3128 383 3136 417
rect 3170 383 3182 417
rect 3128 333 3182 383
rect 3218 333 3287 497
rect 3020 297 3074 309
rect 3235 297 3287 333
rect 3323 485 3377 497
rect 3323 451 3335 485
rect 3369 451 3377 485
rect 3323 417 3377 451
rect 3323 383 3335 417
rect 3369 383 3377 417
rect 3323 349 3377 383
rect 3323 315 3335 349
rect 3369 315 3377 349
rect 3323 297 3377 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 214 82 248 116
rect 338 82 372 116
rect 443 82 477 116
rect 548 82 582 116
rect 672 82 706 116
rect 857 127 891 161
rect 857 59 891 93
rect 1042 82 1076 116
rect 1166 82 1200 116
rect 1271 82 1305 116
rect 1376 82 1410 116
rect 1500 82 1534 116
rect 1685 127 1719 161
rect 1685 59 1719 93
rect 1870 82 1904 116
rect 1994 82 2028 116
rect 2099 82 2133 116
rect 2204 82 2238 116
rect 2328 82 2362 116
rect 2513 127 2547 161
rect 2513 59 2547 93
rect 2698 82 2732 116
rect 2822 82 2856 116
rect 2927 82 2961 116
rect 3032 82 3066 116
rect 3156 82 3190 116
rect 3335 127 3369 161
rect 3335 59 3369 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 234 451 268 485
rect 234 383 268 417
rect 338 445 372 479
rect 338 377 372 411
rect 338 309 372 343
rect 443 445 477 479
rect 443 377 477 411
rect 443 309 477 343
rect 548 445 582 479
rect 548 377 582 411
rect 548 309 582 343
rect 652 451 686 485
rect 652 383 686 417
rect 857 451 891 485
rect 857 383 891 417
rect 857 315 891 349
rect 1062 451 1096 485
rect 1062 383 1096 417
rect 1166 445 1200 479
rect 1166 377 1200 411
rect 1166 309 1200 343
rect 1271 445 1305 479
rect 1271 377 1305 411
rect 1271 309 1305 343
rect 1376 445 1410 479
rect 1376 377 1410 411
rect 1376 309 1410 343
rect 1480 451 1514 485
rect 1480 383 1514 417
rect 1685 451 1719 485
rect 1685 383 1719 417
rect 1685 315 1719 349
rect 1890 451 1924 485
rect 1890 383 1924 417
rect 1994 445 2028 479
rect 1994 377 2028 411
rect 1994 309 2028 343
rect 2099 445 2133 479
rect 2099 377 2133 411
rect 2099 309 2133 343
rect 2204 445 2238 479
rect 2204 377 2238 411
rect 2204 309 2238 343
rect 2308 451 2342 485
rect 2308 383 2342 417
rect 2513 451 2547 485
rect 2513 383 2547 417
rect 2513 315 2547 349
rect 2718 451 2752 485
rect 2718 383 2752 417
rect 2822 445 2856 479
rect 2822 377 2856 411
rect 2822 309 2856 343
rect 2927 445 2961 479
rect 2927 377 2961 411
rect 2927 309 2961 343
rect 3032 445 3066 479
rect 3032 377 3066 411
rect 3032 309 3066 343
rect 3136 451 3170 485
rect 3136 383 3170 417
rect 3335 451 3369 485
rect 3335 383 3369 417
rect 3335 315 3369 349
<< poly >>
rect 81 497 117 523
rect 186 497 222 524
rect 384 497 420 523
rect 500 497 536 523
rect 698 497 734 524
rect 803 497 839 523
rect 909 497 945 523
rect 1014 497 1050 524
rect 1212 497 1248 523
rect 1328 497 1364 523
rect 1526 497 1562 524
rect 1631 497 1667 523
rect 1737 497 1773 523
rect 1842 497 1878 524
rect 2040 497 2076 523
rect 2156 497 2192 523
rect 2354 497 2390 524
rect 2459 497 2495 523
rect 2565 497 2601 523
rect 2670 497 2706 524
rect 2868 497 2904 523
rect 2984 497 3020 523
rect 3182 497 3218 524
rect 3287 497 3323 523
rect 81 282 117 297
rect 186 295 222 333
rect 184 285 298 295
rect 79 265 119 282
rect 184 265 248 285
rect 73 249 127 265
rect 73 215 83 249
rect 117 215 127 249
rect 232 251 248 265
rect 282 251 298 285
rect 384 282 420 297
rect 500 282 536 297
rect 698 295 734 333
rect 622 285 736 295
rect 232 241 298 251
rect 382 239 422 282
rect 73 199 127 215
rect 368 223 422 239
rect 79 177 109 199
rect 368 196 378 223
rect 174 189 378 196
rect 412 189 422 223
rect 174 173 422 189
rect 498 239 538 282
rect 622 251 638 285
rect 672 265 736 285
rect 803 282 839 297
rect 909 282 945 297
rect 1014 295 1050 333
rect 1012 285 1126 295
rect 801 265 841 282
rect 907 265 947 282
rect 1012 265 1076 285
rect 672 251 688 265
rect 622 241 688 251
rect 793 249 847 265
rect 498 223 552 239
rect 498 189 508 223
rect 542 196 552 223
rect 793 215 803 249
rect 837 215 847 249
rect 793 199 847 215
rect 901 249 955 265
rect 901 215 911 249
rect 945 215 955 249
rect 1060 251 1076 265
rect 1110 251 1126 285
rect 1212 282 1248 297
rect 1328 282 1364 297
rect 1526 295 1562 333
rect 1450 285 1564 295
rect 1060 241 1126 251
rect 1210 239 1250 282
rect 901 199 955 215
rect 1196 223 1250 239
rect 542 189 746 196
rect 498 173 746 189
rect 811 177 841 199
rect 907 177 937 199
rect 1196 196 1206 223
rect 1002 189 1206 196
rect 1240 189 1250 223
rect 174 166 417 173
rect 174 151 204 166
rect 387 151 417 166
rect 503 166 746 173
rect 503 151 533 166
rect 716 151 746 166
rect 1002 173 1250 189
rect 1326 239 1366 282
rect 1450 251 1466 285
rect 1500 265 1564 285
rect 1631 282 1667 297
rect 1737 282 1773 297
rect 1842 295 1878 333
rect 1840 285 1954 295
rect 1629 265 1669 282
rect 1735 265 1775 282
rect 1840 265 1904 285
rect 1500 251 1516 265
rect 1450 241 1516 251
rect 1621 249 1675 265
rect 1326 223 1380 239
rect 1326 189 1336 223
rect 1370 196 1380 223
rect 1621 215 1631 249
rect 1665 215 1675 249
rect 1621 199 1675 215
rect 1729 249 1783 265
rect 1729 215 1739 249
rect 1773 215 1783 249
rect 1888 251 1904 265
rect 1938 251 1954 285
rect 2040 282 2076 297
rect 2156 282 2192 297
rect 2354 295 2390 333
rect 2278 285 2392 295
rect 1888 241 1954 251
rect 2038 239 2078 282
rect 1729 199 1783 215
rect 2024 223 2078 239
rect 1370 189 1574 196
rect 1326 173 1574 189
rect 1639 177 1669 199
rect 1735 177 1765 199
rect 2024 196 2034 223
rect 1830 189 2034 196
rect 2068 189 2078 223
rect 1002 166 1245 173
rect 1002 151 1032 166
rect 1215 151 1245 166
rect 1331 166 1574 173
rect 1331 151 1361 166
rect 1544 151 1574 166
rect 1830 173 2078 189
rect 2154 239 2194 282
rect 2278 251 2294 285
rect 2328 265 2392 285
rect 2459 282 2495 297
rect 2565 282 2601 297
rect 2670 295 2706 333
rect 2668 285 2782 295
rect 2457 265 2497 282
rect 2563 265 2603 282
rect 2668 265 2732 285
rect 2328 251 2344 265
rect 2278 241 2344 251
rect 2449 249 2503 265
rect 2154 223 2208 239
rect 2154 189 2164 223
rect 2198 196 2208 223
rect 2449 215 2459 249
rect 2493 215 2503 249
rect 2449 199 2503 215
rect 2557 249 2611 265
rect 2557 215 2567 249
rect 2601 215 2611 249
rect 2716 251 2732 265
rect 2766 251 2782 285
rect 2868 282 2904 297
rect 2984 282 3020 297
rect 3182 295 3218 333
rect 3106 285 3220 295
rect 2716 241 2782 251
rect 2866 239 2906 282
rect 2557 199 2611 215
rect 2852 223 2906 239
rect 2198 189 2402 196
rect 2154 173 2402 189
rect 2467 177 2497 199
rect 2563 177 2593 199
rect 2852 196 2862 223
rect 2658 189 2862 196
rect 2896 189 2906 223
rect 1830 166 2073 173
rect 1830 151 1860 166
rect 2043 151 2073 166
rect 2159 166 2402 173
rect 2159 151 2189 166
rect 2372 151 2402 166
rect 2658 173 2906 189
rect 2982 239 3022 282
rect 3106 251 3122 285
rect 3156 265 3220 285
rect 3287 282 3323 297
rect 3285 265 3325 282
rect 3156 251 3172 265
rect 3106 241 3172 251
rect 3277 249 3331 265
rect 2982 223 3036 239
rect 2982 189 2992 223
rect 3026 196 3036 223
rect 3277 215 3287 249
rect 3321 215 3331 249
rect 3277 199 3331 215
rect 3026 189 3230 196
rect 2982 173 3230 189
rect 3295 177 3325 199
rect 2658 166 2901 173
rect 2658 151 2688 166
rect 2871 151 2901 166
rect 2987 166 3230 173
rect 2987 151 3017 166
rect 3200 151 3230 166
rect 79 21 109 47
rect 174 21 204 47
rect 387 21 417 47
rect 503 21 533 47
rect 716 21 746 47
rect 811 21 841 47
rect 907 21 937 47
rect 1002 21 1032 47
rect 1215 21 1245 47
rect 1331 21 1361 47
rect 1544 21 1574 47
rect 1639 21 1669 47
rect 1735 21 1765 47
rect 1830 21 1860 47
rect 2043 21 2073 47
rect 2159 21 2189 47
rect 2372 21 2402 47
rect 2467 21 2497 47
rect 2563 21 2593 47
rect 2658 21 2688 47
rect 2871 21 2901 47
rect 2987 21 3017 47
rect 3200 21 3230 47
rect 3295 21 3325 47
<< polycont >>
rect 83 215 117 249
rect 248 251 282 285
rect 378 189 412 223
rect 638 251 672 285
rect 508 189 542 223
rect 803 215 837 249
rect 911 215 945 249
rect 1076 251 1110 285
rect 1206 189 1240 223
rect 1466 251 1500 285
rect 1336 189 1370 223
rect 1631 215 1665 249
rect 1739 215 1773 249
rect 1904 251 1938 285
rect 2034 189 2068 223
rect 2294 251 2328 285
rect 2164 189 2198 223
rect 2459 215 2493 249
rect 2567 215 2601 249
rect 2732 251 2766 285
rect 2862 189 2896 223
rect 3122 251 3156 285
rect 2992 189 3026 223
rect 3287 215 3321 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3404 561
rect 19 485 85 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 218 485 284 493
rect 218 451 234 485
rect 268 451 284 485
rect 218 417 284 451
rect 218 397 234 417
rect 19 349 85 383
rect 19 315 35 349
rect 69 315 85 349
rect 19 299 85 315
rect 180 391 234 397
rect 180 357 213 391
rect 268 383 284 417
rect 247 361 284 383
rect 322 479 388 493
rect 322 445 338 479
rect 372 445 388 479
rect 322 411 388 445
rect 322 377 338 411
rect 372 377 388 411
rect 247 357 259 361
rect 180 351 259 357
rect 67 249 146 265
rect 67 215 83 249
rect 117 215 146 249
rect 67 211 146 215
rect 26 161 78 177
rect 26 127 35 161
rect 69 127 78 161
rect 26 93 78 127
rect 26 59 35 93
rect 69 59 78 93
rect 112 125 146 211
rect 180 201 214 351
rect 322 343 388 377
rect 322 327 338 343
rect 292 309 338 327
rect 372 309 388 343
rect 292 301 388 309
rect 248 293 388 301
rect 427 479 493 527
rect 427 445 443 479
rect 477 445 493 479
rect 427 411 493 445
rect 427 377 443 411
rect 477 377 493 411
rect 427 343 493 377
rect 427 309 443 343
rect 477 309 493 343
rect 427 293 493 309
rect 532 479 598 493
rect 532 445 548 479
rect 582 445 598 479
rect 532 411 598 445
rect 532 377 548 411
rect 582 377 598 411
rect 532 343 598 377
rect 636 485 702 493
rect 636 451 652 485
rect 686 451 702 485
rect 636 417 702 451
rect 636 383 652 417
rect 686 397 702 417
rect 835 485 913 527
rect 835 451 857 485
rect 891 451 913 485
rect 835 417 913 451
rect 686 391 740 397
rect 636 361 673 383
rect 661 357 673 361
rect 707 357 740 391
rect 661 351 740 357
rect 532 309 548 343
rect 582 327 598 343
rect 582 309 628 327
rect 532 301 628 309
rect 532 293 672 301
rect 248 285 326 293
rect 282 251 326 285
rect 594 285 672 293
rect 248 235 326 251
rect 180 167 258 201
rect 112 79 167 125
rect 209 116 258 167
rect 292 151 326 235
rect 361 223 441 259
rect 361 189 378 223
rect 412 189 441 223
rect 479 223 559 259
rect 479 189 508 223
rect 542 189 559 223
rect 594 251 638 285
rect 594 235 672 251
rect 594 151 628 235
rect 706 201 740 351
rect 835 383 857 417
rect 891 383 913 417
rect 1046 485 1112 493
rect 1046 451 1062 485
rect 1096 451 1112 485
rect 1046 417 1112 451
rect 1046 397 1062 417
rect 835 349 913 383
rect 835 315 857 349
rect 891 315 913 349
rect 835 299 913 315
rect 1008 391 1062 397
rect 1008 357 1041 391
rect 1096 383 1112 417
rect 1075 361 1112 383
rect 1150 479 1216 493
rect 1150 445 1166 479
rect 1200 445 1216 479
rect 1150 411 1216 445
rect 1150 377 1166 411
rect 1200 377 1216 411
rect 1075 357 1087 361
rect 1008 351 1087 357
rect 292 117 380 151
rect 209 82 214 116
rect 248 82 258 116
rect 209 66 258 82
rect 330 116 380 117
rect 330 82 338 116
rect 372 82 380 116
rect 330 66 380 82
rect 427 116 493 132
rect 427 82 443 116
rect 477 82 493 116
rect 26 17 78 59
rect 427 17 493 82
rect 540 117 628 151
rect 662 167 740 201
rect 774 249 853 265
rect 774 215 803 249
rect 837 215 853 249
rect 774 211 853 215
rect 895 249 974 265
rect 895 215 911 249
rect 945 215 974 249
rect 895 211 974 215
rect 540 116 590 117
rect 540 82 548 116
rect 582 82 590 116
rect 540 66 590 82
rect 662 116 711 167
rect 774 125 808 211
rect 662 82 672 116
rect 706 82 711 116
rect 662 66 711 82
rect 753 79 808 125
rect 842 161 906 177
rect 842 127 857 161
rect 891 127 906 161
rect 842 93 906 127
rect 842 59 857 93
rect 891 59 906 93
rect 940 125 974 211
rect 1008 201 1042 351
rect 1150 343 1216 377
rect 1150 327 1166 343
rect 1120 309 1166 327
rect 1200 309 1216 343
rect 1120 301 1216 309
rect 1076 293 1216 301
rect 1255 479 1321 527
rect 1255 445 1271 479
rect 1305 445 1321 479
rect 1255 411 1321 445
rect 1255 377 1271 411
rect 1305 377 1321 411
rect 1255 343 1321 377
rect 1255 309 1271 343
rect 1305 309 1321 343
rect 1255 293 1321 309
rect 1360 479 1426 493
rect 1360 445 1376 479
rect 1410 445 1426 479
rect 1360 411 1426 445
rect 1360 377 1376 411
rect 1410 377 1426 411
rect 1360 343 1426 377
rect 1464 485 1530 493
rect 1464 451 1480 485
rect 1514 451 1530 485
rect 1464 417 1530 451
rect 1464 383 1480 417
rect 1514 397 1530 417
rect 1663 485 1741 527
rect 1663 451 1685 485
rect 1719 451 1741 485
rect 1663 417 1741 451
rect 1514 391 1568 397
rect 1464 361 1501 383
rect 1489 357 1501 361
rect 1535 357 1568 391
rect 1489 351 1568 357
rect 1360 309 1376 343
rect 1410 327 1426 343
rect 1410 309 1456 327
rect 1360 301 1456 309
rect 1360 293 1500 301
rect 1076 285 1154 293
rect 1110 251 1154 285
rect 1422 285 1500 293
rect 1076 235 1154 251
rect 1008 167 1086 201
rect 940 79 995 125
rect 1037 116 1086 167
rect 1120 151 1154 235
rect 1189 223 1269 259
rect 1189 189 1206 223
rect 1240 189 1269 223
rect 1307 223 1387 259
rect 1307 189 1336 223
rect 1370 189 1387 223
rect 1422 251 1466 285
rect 1422 235 1500 251
rect 1422 151 1456 235
rect 1534 201 1568 351
rect 1663 383 1685 417
rect 1719 383 1741 417
rect 1874 485 1940 493
rect 1874 451 1890 485
rect 1924 451 1940 485
rect 1874 417 1940 451
rect 1874 397 1890 417
rect 1663 349 1741 383
rect 1663 315 1685 349
rect 1719 315 1741 349
rect 1663 299 1741 315
rect 1836 391 1890 397
rect 1836 357 1869 391
rect 1924 383 1940 417
rect 1903 361 1940 383
rect 1978 479 2044 493
rect 1978 445 1994 479
rect 2028 445 2044 479
rect 1978 411 2044 445
rect 1978 377 1994 411
rect 2028 377 2044 411
rect 1903 357 1915 361
rect 1836 351 1915 357
rect 1120 117 1208 151
rect 1037 82 1042 116
rect 1076 82 1086 116
rect 1037 66 1086 82
rect 1158 116 1208 117
rect 1158 82 1166 116
rect 1200 82 1208 116
rect 1158 66 1208 82
rect 1255 116 1321 132
rect 1255 82 1271 116
rect 1305 82 1321 116
rect 842 17 906 59
rect 1255 17 1321 82
rect 1368 117 1456 151
rect 1490 167 1568 201
rect 1602 249 1681 265
rect 1602 215 1631 249
rect 1665 215 1681 249
rect 1602 211 1681 215
rect 1723 249 1802 265
rect 1723 215 1739 249
rect 1773 215 1802 249
rect 1723 211 1802 215
rect 1368 116 1418 117
rect 1368 82 1376 116
rect 1410 82 1418 116
rect 1368 66 1418 82
rect 1490 116 1539 167
rect 1602 125 1636 211
rect 1490 82 1500 116
rect 1534 82 1539 116
rect 1490 66 1539 82
rect 1581 79 1636 125
rect 1670 161 1734 177
rect 1670 127 1685 161
rect 1719 127 1734 161
rect 1670 93 1734 127
rect 1670 59 1685 93
rect 1719 59 1734 93
rect 1768 125 1802 211
rect 1836 201 1870 351
rect 1978 343 2044 377
rect 1978 327 1994 343
rect 1948 309 1994 327
rect 2028 309 2044 343
rect 1948 301 2044 309
rect 1904 293 2044 301
rect 2083 479 2149 527
rect 2083 445 2099 479
rect 2133 445 2149 479
rect 2083 411 2149 445
rect 2083 377 2099 411
rect 2133 377 2149 411
rect 2083 343 2149 377
rect 2083 309 2099 343
rect 2133 309 2149 343
rect 2083 293 2149 309
rect 2188 479 2254 493
rect 2188 445 2204 479
rect 2238 445 2254 479
rect 2188 411 2254 445
rect 2188 377 2204 411
rect 2238 377 2254 411
rect 2188 343 2254 377
rect 2292 485 2358 493
rect 2292 451 2308 485
rect 2342 451 2358 485
rect 2292 417 2358 451
rect 2292 383 2308 417
rect 2342 397 2358 417
rect 2491 485 2569 527
rect 2491 451 2513 485
rect 2547 451 2569 485
rect 2491 417 2569 451
rect 2342 391 2396 397
rect 2292 361 2329 383
rect 2317 357 2329 361
rect 2363 357 2396 391
rect 2317 351 2396 357
rect 2188 309 2204 343
rect 2238 327 2254 343
rect 2238 309 2284 327
rect 2188 301 2284 309
rect 2188 293 2328 301
rect 1904 285 1982 293
rect 1938 251 1982 285
rect 2250 285 2328 293
rect 1904 235 1982 251
rect 1836 167 1914 201
rect 1768 79 1823 125
rect 1865 116 1914 167
rect 1948 151 1982 235
rect 2017 223 2097 259
rect 2017 189 2034 223
rect 2068 189 2097 223
rect 2135 223 2215 259
rect 2135 189 2164 223
rect 2198 189 2215 223
rect 2250 251 2294 285
rect 2250 235 2328 251
rect 2250 151 2284 235
rect 2362 201 2396 351
rect 2491 383 2513 417
rect 2547 383 2569 417
rect 2702 485 2768 493
rect 2702 451 2718 485
rect 2752 451 2768 485
rect 2702 417 2768 451
rect 2702 397 2718 417
rect 2491 349 2569 383
rect 2491 315 2513 349
rect 2547 315 2569 349
rect 2491 299 2569 315
rect 2664 391 2718 397
rect 2664 357 2697 391
rect 2752 383 2768 417
rect 2731 361 2768 383
rect 2806 479 2872 493
rect 2806 445 2822 479
rect 2856 445 2872 479
rect 2806 411 2872 445
rect 2806 377 2822 411
rect 2856 377 2872 411
rect 2731 357 2743 361
rect 2664 351 2743 357
rect 1948 117 2036 151
rect 1865 82 1870 116
rect 1904 82 1914 116
rect 1865 66 1914 82
rect 1986 116 2036 117
rect 1986 82 1994 116
rect 2028 82 2036 116
rect 1986 66 2036 82
rect 2083 116 2149 132
rect 2083 82 2099 116
rect 2133 82 2149 116
rect 1670 17 1734 59
rect 2083 17 2149 82
rect 2196 117 2284 151
rect 2318 167 2396 201
rect 2430 249 2509 265
rect 2430 215 2459 249
rect 2493 215 2509 249
rect 2430 211 2509 215
rect 2551 249 2630 265
rect 2551 215 2567 249
rect 2601 215 2630 249
rect 2551 211 2630 215
rect 2196 116 2246 117
rect 2196 82 2204 116
rect 2238 82 2246 116
rect 2196 66 2246 82
rect 2318 116 2367 167
rect 2430 125 2464 211
rect 2318 82 2328 116
rect 2362 82 2367 116
rect 2318 66 2367 82
rect 2409 79 2464 125
rect 2498 161 2562 177
rect 2498 127 2513 161
rect 2547 127 2562 161
rect 2498 93 2562 127
rect 2498 59 2513 93
rect 2547 59 2562 93
rect 2596 125 2630 211
rect 2664 201 2698 351
rect 2806 343 2872 377
rect 2806 327 2822 343
rect 2776 309 2822 327
rect 2856 309 2872 343
rect 2776 301 2872 309
rect 2732 293 2872 301
rect 2911 479 2977 527
rect 2911 445 2927 479
rect 2961 445 2977 479
rect 2911 411 2977 445
rect 2911 377 2927 411
rect 2961 377 2977 411
rect 2911 343 2977 377
rect 2911 309 2927 343
rect 2961 309 2977 343
rect 2911 293 2977 309
rect 3016 479 3082 493
rect 3016 445 3032 479
rect 3066 445 3082 479
rect 3016 411 3082 445
rect 3016 377 3032 411
rect 3066 377 3082 411
rect 3016 343 3082 377
rect 3120 485 3186 493
rect 3120 451 3136 485
rect 3170 451 3186 485
rect 3120 417 3186 451
rect 3120 383 3136 417
rect 3170 397 3186 417
rect 3319 485 3385 527
rect 3319 451 3335 485
rect 3369 451 3385 485
rect 3319 417 3385 451
rect 3170 391 3224 397
rect 3120 361 3157 383
rect 3145 357 3157 361
rect 3191 357 3224 391
rect 3145 351 3224 357
rect 3016 309 3032 343
rect 3066 327 3082 343
rect 3066 309 3112 327
rect 3016 301 3112 309
rect 3016 293 3156 301
rect 2732 285 2810 293
rect 2766 251 2810 285
rect 3078 285 3156 293
rect 2732 235 2810 251
rect 2664 167 2742 201
rect 2596 79 2651 125
rect 2693 116 2742 167
rect 2776 151 2810 235
rect 2845 223 2925 259
rect 2845 189 2862 223
rect 2896 189 2925 223
rect 2963 223 3043 259
rect 2963 189 2992 223
rect 3026 189 3043 223
rect 3078 251 3122 285
rect 3078 235 3156 251
rect 3078 151 3112 235
rect 3190 201 3224 351
rect 3319 383 3335 417
rect 3369 383 3385 417
rect 3319 349 3385 383
rect 3319 315 3335 349
rect 3369 315 3385 349
rect 3319 299 3385 315
rect 2776 117 2864 151
rect 2693 82 2698 116
rect 2732 82 2742 116
rect 2693 66 2742 82
rect 2814 116 2864 117
rect 2814 82 2822 116
rect 2856 82 2864 116
rect 2814 66 2864 82
rect 2911 116 2977 132
rect 2911 82 2927 116
rect 2961 82 2977 116
rect 2498 17 2562 59
rect 2911 17 2977 82
rect 3024 117 3112 151
rect 3146 167 3224 201
rect 3258 249 3337 265
rect 3258 215 3287 249
rect 3321 215 3337 249
rect 3258 211 3337 215
rect 3024 116 3074 117
rect 3024 82 3032 116
rect 3066 82 3074 116
rect 3024 66 3074 82
rect 3146 116 3195 167
rect 3258 125 3292 211
rect 3146 82 3156 116
rect 3190 82 3195 116
rect 3146 66 3195 82
rect 3237 79 3292 125
rect 3326 161 3378 177
rect 3326 127 3335 161
rect 3369 127 3378 161
rect 3326 93 3378 127
rect 3326 59 3335 93
rect 3369 59 3378 93
rect 3326 17 3378 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3404 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 213 383 234 391
rect 234 383 247 391
rect 213 357 247 383
rect 673 383 686 391
rect 686 383 707 391
rect 673 357 707 383
rect 1041 383 1062 391
rect 1062 383 1075 391
rect 1041 357 1075 383
rect 1501 383 1514 391
rect 1514 383 1535 391
rect 1501 357 1535 383
rect 1869 383 1890 391
rect 1890 383 1903 391
rect 1869 357 1903 383
rect 2329 383 2342 391
rect 2342 383 2363 391
rect 2329 357 2363 383
rect 2697 383 2718 391
rect 2718 383 2731 391
rect 2697 357 2731 383
rect 3157 383 3170 391
rect 3170 383 3191 391
rect 3157 357 3191 383
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
<< metal1 >>
rect 0 561 3404 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3404 561
rect 0 496 3404 527
rect 201 391 259 397
rect 201 357 213 391
rect 247 388 259 391
rect 661 391 719 397
rect 661 388 673 391
rect 247 360 673 388
rect 247 357 259 360
rect 201 351 259 357
rect 661 357 673 360
rect 707 388 719 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 707 360 1041 388
rect 707 357 719 360
rect 661 351 719 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1489 391 1547 397
rect 1489 388 1501 391
rect 1075 360 1501 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1489 357 1501 360
rect 1535 388 1547 391
rect 1857 391 1915 397
rect 1857 388 1869 391
rect 1535 360 1869 388
rect 1535 357 1547 360
rect 1489 351 1547 357
rect 1857 357 1869 360
rect 1903 388 1915 391
rect 2317 391 2375 397
rect 2317 388 2329 391
rect 1903 360 2329 388
rect 1903 357 1915 360
rect 1857 351 1915 357
rect 2317 357 2329 360
rect 2363 388 2375 391
rect 2685 391 2743 397
rect 2685 388 2697 391
rect 2363 360 2697 388
rect 2363 357 2375 360
rect 2317 351 2375 357
rect 2685 357 2697 360
rect 2731 388 2743 391
rect 3145 391 3203 397
rect 3145 388 3157 391
rect 2731 360 3157 388
rect 2731 357 2743 360
rect 2685 351 2743 357
rect 3145 357 3157 360
rect 3191 357 3203 391
rect 3145 351 3203 357
rect 0 17 3404 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3404 17
rect 0 -48 3404 -17
<< labels >>
rlabel comment s 0 0 0 0 4 muxb8to1_1
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 17 nsew ground bidirectional
flabel metal1 s 213 357 247 391 0 FreeSans 200 0 0 0 Z
port 21 nsew signal output
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 20 nsew power bidirectional
flabel metal1 s 3157 357 3191 391 0 FreeSans 200 180 0 0 Z
port 21 nsew signal output
flabel metal1 s 3341 527 3375 561 0 FreeSans 200 180 0 0 VPWR
port 20 nsew power bidirectional
flabel metal1 s 3341 -17 3375 17 0 FreeSans 200 180 0 0 VGND
port 17 nsew ground bidirectional
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 230 374 230 374 0 FreeSans 200 0 0 0 Z
flabel metal1 s 2697 357 2731 391 0 FreeSans 200 0 0 0 Z
port 21 nsew
flabel metal1 s 2513 527 2547 561 0 FreeSans 200 0 0 0 VPWR
port 20 nsew
flabel metal1 s 2513 -17 2547 17 0 FreeSans 200 0 0 0 VGND
port 17 nsew
flabel metal1 s 2329 357 2363 391 0 FreeSans 200 180 0 0 Z
port 21 nsew
flabel metal1 s 2530 544 2530 544 0 FreeSans 200 180 0 0 VPWR
flabel metal1 s 2530 0 2530 0 0 FreeSans 200 180 0 0 VGND
flabel metal1 s 1501 357 1535 391 0 FreeSans 200 180 0 0 Z
port 21 nsew
flabel metal1 s 1685 527 1719 561 0 FreeSans 200 180 0 0 VPWR
port 20 nsew
flabel metal1 s 1685 -17 1719 17 0 FreeSans 200 180 0 0 VGND
port 17 nsew
flabel metal1 s 1869 357 1903 391 0 FreeSans 200 0 0 0 Z
port 21 nsew
flabel metal1 s 1702 544 1702 544 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 1702 0 1702 0 0 FreeSans 200 0 0 0 VGND
flabel metal1 s 673 357 707 391 0 FreeSans 200 180 0 0 Z
port 21 nsew
flabel metal1 s 857 527 891 561 0 FreeSans 200 180 0 0 VPWR
port 20 nsew
flabel metal1 s 857 -17 891 17 0 FreeSans 200 180 0 0 VGND
port 17 nsew
flabel metal1 s 1041 357 1075 391 0 FreeSans 200 0 0 0 Z
port 21 nsew
flabel metal1 s 874 544 874 544 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 874 0 874 0 0 FreeSans 200 0 0 0 VGND
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 18 nsew ground bidirectional
flabel pwell s 3341 -17 3375 17 0 FreeSans 200 180 0 0 VNB
port 18 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel pwell s 2513 -17 2547 17 0 FreeSans 200 0 0 0 VNB
port 18 nsew
flabel pwell s 2530 0 2530 0 0 FreeSans 200 180 0 0 VNB
flabel pwell s 1685 -17 1719 17 0 FreeSans 200 180 0 0 VNB
port 18 nsew
flabel pwell s 1702 0 1702 0 0 FreeSans 200 0 0 0 VNB
flabel pwell s 857 -17 891 17 0 FreeSans 200 180 0 0 VNB
port 18 nsew
flabel pwell s 874 0 874 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 19 nsew power bidirectional
flabel nwell s 3341 527 3375 561 0 FreeSans 200 180 0 0 VPB
port 19 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel nwell s 2513 527 2547 561 0 FreeSans 200 0 0 0 VPB
port 19 nsew
flabel nwell s 2530 544 2530 544 0 FreeSans 200 180 0 0 VPB
flabel nwell s 1685 527 1719 561 0 FreeSans 200 180 0 0 VPB
port 19 nsew
flabel nwell s 1702 544 1702 544 0 FreeSans 200 0 0 0 VPB
flabel nwell s 857 527 891 561 0 FreeSans 200 180 0 0 VPB
port 19 nsew
flabel nwell s 874 544 874 544 0 FreeSans 200 0 0 0 VPB
flabel locali s 121 85 155 119 0 FreeSans 200 0 0 0 D[0]
port 8 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 S[0]
port 16 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 S[1]
port 15 nsew signal input
flabel locali s 765 85 799 119 0 FreeSans 200 0 0 0 D[1]
port 7 nsew signal input
flabel locali s 949 85 983 119 0 FreeSans 200 0 0 0 D[2]
port 6 nsew signal input
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 S[2]
port 14 nsew signal input
flabel locali s 1317 221 1351 255 0 FreeSans 200 0 0 0 S[3]
port 13 nsew signal input
flabel locali s 1777 85 1811 119 0 FreeSans 200 0 0 0 D[4]
port 4 nsew signal input
flabel locali s 2053 221 2087 255 0 FreeSans 200 0 0 0 S[4]
port 12 nsew signal input
flabel locali s 2145 221 2179 255 0 FreeSans 200 0 0 0 S[5]
port 11 nsew signal input
flabel locali s 2421 85 2455 119 0 FreeSans 200 0 0 0 D[5]
port 3 nsew signal input
flabel locali s 2605 85 2639 119 0 FreeSans 200 0 0 0 D[6]
port 2 nsew signal input
flabel locali s 2881 221 2915 255 0 FreeSans 200 0 0 0 S[6]
port 10 nsew signal input
flabel locali s 2973 221 3007 255 0 FreeSans 200 0 0 0 S[7]
port 9 nsew signal input
flabel locali s 3249 85 3283 119 0 FreeSans 200 0 0 0 D[7]
port 1 nsew signal input
flabel locali s 1593 85 1627 119 0 FreeSans 200 0 0 0 D[3]
port 5 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 3404 544
string GDS_END 3056860
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 3009326
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
