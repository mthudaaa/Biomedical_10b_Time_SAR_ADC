magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 215 21 1581 157
rect 30 -17 64 17
<< scnmos >>
rect 371 47 401 131
rect 455 47 485 131
rect 559 47 589 131
rect 643 47 673 131
rect 747 47 777 131
rect 831 47 861 131
rect 935 47 965 131
rect 1019 47 1049 131
rect 1123 47 1153 131
rect 1207 47 1237 131
rect 1311 47 1341 131
rect 1395 47 1425 131
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
rect 1209 297 1245 497
rect 1303 297 1339 497
rect 1397 297 1433 497
rect 1491 297 1527 497
rect 1585 297 1621 497
rect 1679 297 1715 497
<< ndiff >>
rect 241 97 371 131
rect 241 63 249 97
rect 283 63 317 97
rect 351 63 371 97
rect 241 47 371 63
rect 401 106 455 131
rect 401 72 411 106
rect 445 72 455 106
rect 401 47 455 72
rect 485 97 559 131
rect 485 63 505 97
rect 539 63 559 97
rect 485 47 559 63
rect 589 106 643 131
rect 589 72 599 106
rect 633 72 643 106
rect 589 47 643 72
rect 673 97 747 131
rect 673 63 693 97
rect 727 63 747 97
rect 673 47 747 63
rect 777 106 831 131
rect 777 72 787 106
rect 821 72 831 106
rect 777 47 831 72
rect 861 97 935 131
rect 861 63 881 97
rect 915 63 935 97
rect 861 47 935 63
rect 965 106 1019 131
rect 965 72 975 106
rect 1009 72 1019 106
rect 965 47 1019 72
rect 1049 97 1123 131
rect 1049 63 1069 97
rect 1103 63 1123 97
rect 1049 47 1123 63
rect 1153 106 1207 131
rect 1153 72 1163 106
rect 1197 72 1207 106
rect 1153 47 1207 72
rect 1237 97 1311 131
rect 1237 63 1257 97
rect 1291 63 1311 97
rect 1237 47 1311 63
rect 1341 106 1395 131
rect 1341 72 1351 106
rect 1385 72 1395 106
rect 1341 47 1395 72
rect 1425 97 1555 131
rect 1425 63 1445 97
rect 1479 63 1513 97
rect 1547 63 1555 97
rect 1425 47 1555 63
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 402 81 451
rect 27 368 35 402
rect 69 368 81 402
rect 27 297 81 368
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 341 175 375
rect 117 307 129 341
rect 163 307 175 341
rect 117 297 175 307
rect 211 489 269 497
rect 211 455 223 489
rect 257 455 269 489
rect 211 402 269 455
rect 211 368 223 402
rect 257 368 269 402
rect 211 297 269 368
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 409 363 443
rect 305 375 317 409
rect 351 375 363 409
rect 305 341 363 375
rect 305 307 317 341
rect 351 307 363 341
rect 305 297 363 307
rect 399 489 457 497
rect 399 455 411 489
rect 445 455 457 489
rect 399 402 457 455
rect 399 368 411 402
rect 445 368 457 402
rect 399 297 457 368
rect 493 477 551 497
rect 493 443 505 477
rect 539 443 551 477
rect 493 409 551 443
rect 493 375 505 409
rect 539 375 551 409
rect 493 341 551 375
rect 493 307 505 341
rect 539 307 551 341
rect 493 297 551 307
rect 587 489 645 497
rect 587 455 599 489
rect 633 455 645 489
rect 587 402 645 455
rect 587 368 599 402
rect 633 368 645 402
rect 587 297 645 368
rect 681 477 739 497
rect 681 443 693 477
rect 727 443 739 477
rect 681 409 739 443
rect 681 375 693 409
rect 727 375 739 409
rect 681 341 739 375
rect 681 307 693 341
rect 727 307 739 341
rect 681 297 739 307
rect 775 489 833 497
rect 775 455 787 489
rect 821 455 833 489
rect 775 402 833 455
rect 775 368 787 402
rect 821 368 833 402
rect 775 297 833 368
rect 869 477 927 497
rect 869 443 881 477
rect 915 443 927 477
rect 869 409 927 443
rect 869 375 881 409
rect 915 375 927 409
rect 869 341 927 375
rect 869 307 881 341
rect 915 307 927 341
rect 869 297 927 307
rect 963 489 1021 497
rect 963 455 975 489
rect 1009 455 1021 489
rect 963 402 1021 455
rect 963 368 975 402
rect 1009 368 1021 402
rect 963 297 1021 368
rect 1057 477 1115 497
rect 1057 443 1069 477
rect 1103 443 1115 477
rect 1057 409 1115 443
rect 1057 375 1069 409
rect 1103 375 1115 409
rect 1057 341 1115 375
rect 1057 307 1069 341
rect 1103 307 1115 341
rect 1057 297 1115 307
rect 1151 489 1209 497
rect 1151 455 1163 489
rect 1197 455 1209 489
rect 1151 402 1209 455
rect 1151 368 1163 402
rect 1197 368 1209 402
rect 1151 297 1209 368
rect 1245 477 1303 497
rect 1245 443 1257 477
rect 1291 443 1303 477
rect 1245 409 1303 443
rect 1245 375 1257 409
rect 1291 375 1303 409
rect 1245 341 1303 375
rect 1245 307 1257 341
rect 1291 307 1303 341
rect 1245 297 1303 307
rect 1339 489 1397 497
rect 1339 455 1351 489
rect 1385 455 1397 489
rect 1339 402 1397 455
rect 1339 368 1351 402
rect 1385 368 1397 402
rect 1339 297 1397 368
rect 1433 477 1491 497
rect 1433 443 1445 477
rect 1479 443 1491 477
rect 1433 409 1491 443
rect 1433 375 1445 409
rect 1479 375 1491 409
rect 1433 341 1491 375
rect 1433 307 1445 341
rect 1479 307 1491 341
rect 1433 297 1491 307
rect 1527 489 1585 497
rect 1527 455 1539 489
rect 1573 455 1585 489
rect 1527 402 1585 455
rect 1527 368 1539 402
rect 1573 368 1585 402
rect 1527 297 1585 368
rect 1621 477 1679 497
rect 1621 443 1633 477
rect 1667 443 1679 477
rect 1621 409 1679 443
rect 1621 375 1633 409
rect 1667 375 1679 409
rect 1621 341 1679 375
rect 1621 307 1633 341
rect 1667 307 1679 341
rect 1621 297 1679 307
rect 1715 485 1769 497
rect 1715 451 1727 485
rect 1761 451 1769 485
rect 1715 402 1769 451
rect 1715 368 1727 402
rect 1761 368 1769 402
rect 1715 297 1769 368
<< ndiffc >>
rect 249 63 283 97
rect 317 63 351 97
rect 411 72 445 106
rect 505 63 539 97
rect 599 72 633 106
rect 693 63 727 97
rect 787 72 821 106
rect 881 63 915 97
rect 975 72 1009 106
rect 1069 63 1103 97
rect 1163 72 1197 106
rect 1257 63 1291 97
rect 1351 72 1385 106
rect 1445 63 1479 97
rect 1513 63 1547 97
<< pdiffc >>
rect 35 451 69 485
rect 35 368 69 402
rect 129 443 163 477
rect 129 375 163 409
rect 129 307 163 341
rect 223 455 257 489
rect 223 368 257 402
rect 317 443 351 477
rect 317 375 351 409
rect 317 307 351 341
rect 411 455 445 489
rect 411 368 445 402
rect 505 443 539 477
rect 505 375 539 409
rect 505 307 539 341
rect 599 455 633 489
rect 599 368 633 402
rect 693 443 727 477
rect 693 375 727 409
rect 693 307 727 341
rect 787 455 821 489
rect 787 368 821 402
rect 881 443 915 477
rect 881 375 915 409
rect 881 307 915 341
rect 975 455 1009 489
rect 975 368 1009 402
rect 1069 443 1103 477
rect 1069 375 1103 409
rect 1069 307 1103 341
rect 1163 455 1197 489
rect 1163 368 1197 402
rect 1257 443 1291 477
rect 1257 375 1291 409
rect 1257 307 1291 341
rect 1351 455 1385 489
rect 1351 368 1385 402
rect 1445 443 1479 477
rect 1445 375 1479 409
rect 1445 307 1479 341
rect 1539 455 1573 489
rect 1539 368 1573 402
rect 1633 443 1667 477
rect 1633 375 1667 409
rect 1633 307 1667 341
rect 1727 451 1761 485
rect 1727 368 1761 402
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 1209 497 1245 523
rect 1303 497 1339 523
rect 1397 497 1433 523
rect 1491 497 1527 523
rect 1585 497 1621 523
rect 1679 497 1715 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 1209 282 1245 297
rect 1303 282 1339 297
rect 1397 282 1433 297
rect 1491 282 1527 297
rect 1585 282 1621 297
rect 1679 282 1715 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 831 265 871 282
rect 925 265 965 282
rect 1019 265 1059 282
rect 1113 265 1153 282
rect 1207 265 1247 282
rect 1301 265 1341 282
rect 1395 265 1435 282
rect 1489 265 1529 282
rect 1583 265 1623 282
rect 1677 265 1717 282
rect 79 249 1717 265
rect 79 215 107 249
rect 141 215 175 249
rect 209 215 243 249
rect 277 215 311 249
rect 345 215 379 249
rect 413 215 447 249
rect 481 215 515 249
rect 549 215 583 249
rect 617 215 651 249
rect 685 215 719 249
rect 753 215 787 249
rect 821 215 855 249
rect 889 215 923 249
rect 957 215 991 249
rect 1025 215 1059 249
rect 1093 215 1127 249
rect 1161 215 1195 249
rect 1229 215 1263 249
rect 1297 215 1331 249
rect 1365 215 1399 249
rect 1433 215 1467 249
rect 1501 215 1535 249
rect 1569 215 1717 249
rect 79 199 1717 215
rect 371 131 401 199
rect 455 131 485 199
rect 559 131 589 199
rect 643 131 673 199
rect 747 131 777 199
rect 831 131 861 199
rect 935 131 965 199
rect 1019 131 1049 199
rect 1123 131 1153 199
rect 1207 131 1237 199
rect 1311 131 1341 199
rect 1395 131 1425 199
rect 371 21 401 47
rect 455 21 485 47
rect 559 21 589 47
rect 643 21 673 47
rect 747 21 777 47
rect 831 21 861 47
rect 935 21 965 47
rect 1019 21 1049 47
rect 1123 21 1153 47
rect 1207 21 1237 47
rect 1311 21 1341 47
rect 1395 21 1425 47
<< polycont >>
rect 107 215 141 249
rect 175 215 209 249
rect 243 215 277 249
rect 311 215 345 249
rect 379 215 413 249
rect 447 215 481 249
rect 515 215 549 249
rect 583 215 617 249
rect 651 215 685 249
rect 719 215 753 249
rect 787 215 821 249
rect 855 215 889 249
rect 923 215 957 249
rect 991 215 1025 249
rect 1059 215 1093 249
rect 1127 215 1161 249
rect 1195 215 1229 249
rect 1263 215 1297 249
rect 1331 215 1365 249
rect 1399 215 1433 249
rect 1467 215 1501 249
rect 1535 215 1569 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 19 485 85 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 402 85 451
rect 19 368 35 402
rect 69 368 85 402
rect 19 360 85 368
rect 119 477 173 493
rect 119 443 129 477
rect 163 443 173 477
rect 119 409 173 443
rect 119 375 129 409
rect 163 375 173 409
rect 119 341 173 375
rect 207 489 273 527
rect 207 455 223 489
rect 257 455 273 489
rect 207 402 273 455
rect 207 368 223 402
rect 257 368 273 402
rect 207 360 273 368
rect 307 477 361 493
rect 307 443 317 477
rect 351 443 361 477
rect 307 409 361 443
rect 307 375 317 409
rect 351 375 361 409
rect 119 326 129 341
rect 23 307 129 326
rect 163 326 173 341
rect 307 341 361 375
rect 395 489 461 527
rect 395 455 411 489
rect 445 455 461 489
rect 395 402 461 455
rect 395 368 411 402
rect 445 368 461 402
rect 395 360 461 368
rect 495 477 549 493
rect 495 443 505 477
rect 539 443 549 477
rect 495 409 549 443
rect 495 375 505 409
rect 539 375 549 409
rect 307 326 317 341
rect 163 307 317 326
rect 351 326 361 341
rect 495 341 549 375
rect 583 489 649 527
rect 583 455 599 489
rect 633 455 649 489
rect 583 402 649 455
rect 583 368 599 402
rect 633 368 649 402
rect 583 360 649 368
rect 683 477 737 493
rect 683 443 693 477
rect 727 443 737 477
rect 683 409 737 443
rect 683 375 693 409
rect 727 375 737 409
rect 495 326 505 341
rect 351 307 505 326
rect 539 326 549 341
rect 683 341 737 375
rect 771 489 837 527
rect 771 455 787 489
rect 821 455 837 489
rect 771 402 837 455
rect 771 368 787 402
rect 821 368 837 402
rect 771 360 837 368
rect 871 477 925 493
rect 871 443 881 477
rect 915 443 925 477
rect 871 409 925 443
rect 871 375 881 409
rect 915 375 925 409
rect 683 326 693 341
rect 539 307 693 326
rect 727 326 737 341
rect 871 341 925 375
rect 959 489 1025 527
rect 959 455 975 489
rect 1009 455 1025 489
rect 959 402 1025 455
rect 959 368 975 402
rect 1009 368 1025 402
rect 959 360 1025 368
rect 1059 477 1113 493
rect 1059 443 1069 477
rect 1103 443 1113 477
rect 1059 409 1113 443
rect 1059 375 1069 409
rect 1103 375 1113 409
rect 871 326 881 341
rect 727 307 881 326
rect 915 326 925 341
rect 1059 341 1113 375
rect 1147 489 1213 527
rect 1147 455 1163 489
rect 1197 455 1213 489
rect 1147 402 1213 455
rect 1147 368 1163 402
rect 1197 368 1213 402
rect 1147 360 1213 368
rect 1247 477 1301 493
rect 1247 443 1257 477
rect 1291 443 1301 477
rect 1247 409 1301 443
rect 1247 375 1257 409
rect 1291 375 1301 409
rect 1059 326 1069 341
rect 915 307 1069 326
rect 1103 326 1113 341
rect 1247 341 1301 375
rect 1335 489 1401 527
rect 1335 455 1351 489
rect 1385 455 1401 489
rect 1335 402 1401 455
rect 1335 368 1351 402
rect 1385 368 1401 402
rect 1335 360 1401 368
rect 1435 477 1489 493
rect 1435 443 1445 477
rect 1479 443 1489 477
rect 1435 409 1489 443
rect 1435 375 1445 409
rect 1479 375 1489 409
rect 1247 326 1257 341
rect 1103 307 1257 326
rect 1291 326 1301 341
rect 1435 341 1489 375
rect 1523 489 1589 527
rect 1523 455 1539 489
rect 1573 455 1589 489
rect 1523 402 1589 455
rect 1523 368 1539 402
rect 1573 368 1589 402
rect 1523 360 1589 368
rect 1623 477 1677 493
rect 1623 443 1633 477
rect 1667 443 1677 477
rect 1623 409 1677 443
rect 1623 375 1633 409
rect 1667 375 1677 409
rect 1435 326 1445 341
rect 1291 307 1445 326
rect 1479 326 1489 341
rect 1623 341 1677 375
rect 1711 485 1777 527
rect 1711 451 1727 485
rect 1761 451 1777 485
rect 1711 402 1777 451
rect 1711 368 1727 402
rect 1761 368 1777 402
rect 1711 360 1777 368
rect 1623 326 1633 341
rect 1479 307 1633 326
rect 1667 326 1677 341
rect 1667 307 1731 326
rect 23 292 1731 307
rect 23 173 57 292
rect 91 249 1585 258
rect 91 215 107 249
rect 141 215 175 249
rect 209 215 243 249
rect 277 215 311 249
rect 345 215 379 249
rect 413 215 447 249
rect 481 215 515 249
rect 549 215 583 249
rect 617 215 651 249
rect 685 215 719 249
rect 753 215 787 249
rect 821 215 855 249
rect 889 215 923 249
rect 957 215 991 249
rect 1025 215 1059 249
rect 1093 215 1127 249
rect 1161 215 1195 249
rect 1229 215 1263 249
rect 1297 215 1331 249
rect 1365 215 1399 249
rect 1433 215 1467 249
rect 1501 215 1535 249
rect 1569 215 1585 249
rect 91 207 1585 215
rect 1620 173 1731 292
rect 23 139 1731 173
rect 401 106 455 139
rect 233 97 367 105
rect 233 63 249 97
rect 283 63 317 97
rect 351 63 367 97
rect 233 17 367 63
rect 401 72 411 106
rect 445 72 455 106
rect 589 106 643 139
rect 401 51 455 72
rect 489 97 555 105
rect 489 63 505 97
rect 539 63 555 97
rect 489 17 555 63
rect 589 72 599 106
rect 633 72 643 106
rect 777 106 831 139
rect 589 51 643 72
rect 677 97 743 105
rect 677 63 693 97
rect 727 63 743 97
rect 677 17 743 63
rect 777 72 787 106
rect 821 72 831 106
rect 965 106 1019 139
rect 777 51 831 72
rect 865 97 931 105
rect 865 63 881 97
rect 915 63 931 97
rect 865 17 931 63
rect 965 72 975 106
rect 1009 72 1019 106
rect 1153 106 1207 139
rect 965 51 1019 72
rect 1053 97 1119 105
rect 1053 63 1069 97
rect 1103 63 1119 97
rect 1053 17 1119 63
rect 1153 72 1163 106
rect 1197 72 1207 106
rect 1341 106 1395 139
rect 1153 51 1207 72
rect 1241 97 1307 105
rect 1241 63 1257 97
rect 1291 63 1307 97
rect 1241 17 1307 63
rect 1341 72 1351 106
rect 1385 72 1395 106
rect 1341 51 1395 72
rect 1429 97 1563 105
rect 1429 63 1445 97
rect 1479 63 1513 97
rect 1547 63 1563 97
rect 1429 17 1563 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel locali s 1685 221 1719 255 0 FreeSans 400 0 0 0 Y
port 6 nsew signal output
flabel locali s 857 221 891 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkinv_12
<< properties >>
string FIXED_BBOX 0 0 1840 544
string GDS_END 154940
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 142560
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
