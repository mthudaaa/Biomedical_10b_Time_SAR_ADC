magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 805 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 175 47 205 177
rect 391 47 421 177
rect 470 47 500 177
rect 579 47 609 177
rect 687 47 717 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 383 297 419 497
rect 499 297 535 497
rect 607 297 643 497
rect 689 297 725 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 93 79 131
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 169 175 177
rect 109 135 130 169
rect 164 135 175 169
rect 109 101 175 135
rect 109 67 129 101
rect 163 67 175 101
rect 109 47 175 67
rect 205 89 391 177
rect 205 55 225 89
rect 259 55 294 89
rect 328 55 391 89
rect 205 47 391 55
rect 421 47 470 177
rect 500 157 579 177
rect 500 123 521 157
rect 555 123 579 157
rect 500 89 579 123
rect 500 55 521 89
rect 555 55 579 89
rect 500 47 579 55
rect 609 89 687 177
rect 609 55 637 89
rect 671 55 687 89
rect 609 47 687 55
rect 717 165 779 177
rect 717 131 737 165
rect 771 131 779 165
rect 717 97 779 131
rect 717 63 737 97
rect 771 63 779 97
rect 717 47 779 63
<< pdiff >>
rect 27 484 81 497
rect 27 450 35 484
rect 69 450 81 484
rect 27 416 81 450
rect 27 382 35 416
rect 69 382 81 416
rect 27 348 81 382
rect 27 314 35 348
rect 69 314 81 348
rect 27 297 81 314
rect 117 430 175 497
rect 117 396 129 430
rect 163 396 175 430
rect 117 342 175 396
rect 117 308 129 342
rect 163 308 175 342
rect 117 297 175 308
rect 211 485 265 497
rect 211 451 223 485
rect 257 451 265 485
rect 211 417 265 451
rect 211 383 223 417
rect 257 383 265 417
rect 211 297 265 383
rect 319 485 383 497
rect 319 451 327 485
rect 361 451 383 485
rect 319 417 383 451
rect 319 383 327 417
rect 361 383 383 417
rect 319 297 383 383
rect 419 488 499 497
rect 419 454 444 488
rect 478 454 499 488
rect 419 297 499 454
rect 535 485 607 497
rect 535 451 559 485
rect 593 451 607 485
rect 535 417 607 451
rect 535 383 559 417
rect 593 383 607 417
rect 535 297 607 383
rect 643 297 689 497
rect 725 436 779 497
rect 725 402 737 436
rect 771 402 779 436
rect 725 368 779 402
rect 725 334 737 368
rect 771 334 779 368
rect 725 297 779 334
<< ndiffc >>
rect 35 131 69 165
rect 35 59 69 93
rect 130 135 164 169
rect 129 67 163 101
rect 225 55 259 89
rect 294 55 328 89
rect 521 123 555 157
rect 521 55 555 89
rect 637 55 671 89
rect 737 131 771 165
rect 737 63 771 97
<< pdiffc >>
rect 35 450 69 484
rect 35 382 69 416
rect 35 314 69 348
rect 129 396 163 430
rect 129 308 163 342
rect 223 451 257 485
rect 223 383 257 417
rect 327 451 361 485
rect 327 383 361 417
rect 444 454 478 488
rect 559 451 593 485
rect 559 383 593 417
rect 737 402 771 436
rect 737 334 771 368
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 383 497 419 523
rect 499 497 535 523
rect 607 497 643 523
rect 689 497 725 523
rect 81 282 117 297
rect 175 282 211 297
rect 383 282 419 297
rect 499 282 535 297
rect 607 282 643 297
rect 689 282 725 297
rect 79 265 119 282
rect 173 265 213 282
rect 381 265 421 282
rect 497 265 537 282
rect 605 265 645 282
rect 79 249 264 265
rect 79 215 220 249
rect 254 215 264 249
rect 79 200 264 215
rect 79 177 109 200
rect 175 199 264 200
rect 322 249 421 265
rect 322 215 332 249
rect 366 215 421 249
rect 322 199 421 215
rect 175 177 205 199
rect 391 177 421 199
rect 470 249 537 265
rect 470 215 480 249
rect 514 215 537 249
rect 470 199 537 215
rect 579 249 645 265
rect 579 215 589 249
rect 623 215 645 249
rect 579 199 645 215
rect 687 265 727 282
rect 687 249 741 265
rect 687 215 697 249
rect 731 215 741 249
rect 687 199 741 215
rect 470 177 500 199
rect 579 177 609 199
rect 687 177 717 199
rect 79 21 109 47
rect 175 21 205 47
rect 391 21 421 47
rect 470 21 500 47
rect 579 21 609 47
rect 687 21 717 47
<< polycont >>
rect 220 215 254 249
rect 332 215 366 249
rect 480 215 514 249
rect 589 215 623 249
rect 697 215 731 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 484 77 527
rect 18 450 35 484
rect 69 450 77 484
rect 220 485 271 527
rect 18 416 77 450
rect 18 382 35 416
rect 69 382 77 416
rect 18 348 77 382
rect 18 314 35 348
rect 69 314 77 348
rect 18 298 77 314
rect 121 430 167 467
rect 121 396 129 430
rect 163 396 167 430
rect 121 342 167 396
rect 220 451 223 485
rect 257 451 271 485
rect 220 417 271 451
rect 220 383 223 417
rect 257 383 271 417
rect 220 366 271 383
rect 311 485 387 493
rect 311 451 327 485
rect 361 451 387 485
rect 311 417 387 451
rect 431 488 486 527
rect 431 454 444 488
rect 478 454 486 488
rect 431 438 486 454
rect 543 485 609 493
rect 543 451 559 485
rect 593 451 609 485
rect 311 383 327 417
rect 361 404 387 417
rect 543 417 609 451
rect 543 404 559 417
rect 361 383 559 404
rect 593 383 609 417
rect 311 368 609 383
rect 711 436 787 465
rect 711 402 737 436
rect 771 402 787 436
rect 711 368 787 402
rect 121 308 129 342
rect 163 308 167 342
rect 711 334 737 368
rect 771 334 787 368
rect 711 332 787 334
rect 18 165 77 181
rect 18 131 35 165
rect 69 131 77 165
rect 18 93 77 131
rect 18 59 35 93
rect 69 59 77 93
rect 18 17 77 59
rect 121 169 167 308
rect 121 135 130 169
rect 164 135 167 169
rect 220 298 787 332
rect 220 249 271 298
rect 254 215 271 249
rect 220 175 271 215
rect 305 249 392 255
rect 305 215 332 249
rect 366 215 392 249
rect 305 209 392 215
rect 458 249 539 255
rect 458 215 480 249
rect 514 215 539 249
rect 458 209 539 215
rect 573 249 639 255
rect 573 215 589 249
rect 623 215 639 249
rect 573 209 639 215
rect 673 249 747 255
rect 673 215 697 249
rect 731 215 747 249
rect 673 209 747 215
rect 220 165 787 175
rect 220 157 737 165
rect 220 139 521 157
rect 121 101 167 135
rect 121 67 129 101
rect 163 67 167 101
rect 495 123 521 139
rect 555 139 737 157
rect 555 123 571 139
rect 495 89 571 123
rect 711 131 737 139
rect 771 131 787 165
rect 121 51 167 67
rect 201 55 225 89
rect 259 55 294 89
rect 328 55 354 89
rect 495 55 521 89
rect 555 55 571 89
rect 622 89 677 105
rect 622 55 637 89
rect 671 55 677 89
rect 711 97 787 131
rect 711 63 737 97
rect 771 63 787 97
rect 711 55 787 63
rect 201 17 354 55
rect 622 17 677 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 132 425 166 459 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 305 209 392 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 487 221 521 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 595 221 629 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 700 221 734 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a211o_2
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 29926
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 23234
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
