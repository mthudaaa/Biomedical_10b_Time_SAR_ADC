magic
tech sky130A
magscale 1 2
timestamp 1729608623
<< nwell >>
rect 729 2293 3468 2614
rect 739 1772 907 1777
rect 729 1771 1909 1772
rect 729 1205 3402 1771
rect 2423 362 2612 683
rect 3336 520 3454 683
rect 3329 450 3454 520
rect 3336 362 3454 450
<< psubdiff >>
rect 723 2049 759 2073
rect 723 2015 724 2049
rect 758 2015 759 2049
rect 723 1991 759 2015
rect 704 961 740 985
rect 704 927 705 961
rect 739 927 740 961
rect 704 903 740 927
<< nsubdiff >>
rect 3350 2483 3432 2507
rect 3350 2449 3374 2483
rect 3408 2449 3432 2483
rect 3350 2425 3432 2449
rect 3284 1505 3366 1529
rect 3284 1471 3308 1505
rect 3342 1471 3366 1505
rect 3284 1447 3366 1471
rect 3336 527 3418 551
rect 3336 493 3360 527
rect 3394 493 3418 527
rect 3336 469 3418 493
<< psubdiffcont >>
rect 724 2015 758 2049
rect 705 927 739 961
<< nsubdiffcont >>
rect 3374 2449 3408 2483
rect 3308 1471 3342 1505
rect 3360 493 3394 527
<< locali >>
rect 3350 2483 3432 2507
rect 3350 2449 3374 2483
rect 3408 2449 3432 2483
rect 3350 2425 3432 2449
rect 724 2049 758 2065
rect 758 2015 798 2049
rect 724 1999 758 2015
rect 3284 1505 3366 1529
rect 3284 1471 3308 1505
rect 3342 1471 3366 1505
rect 3284 1447 3366 1471
rect 705 961 739 977
rect 739 927 790 961
rect 3227 927 3317 961
rect 705 911 739 927
rect 3336 527 3418 551
rect 3336 493 3360 527
rect 3394 493 3418 527
rect 3336 469 3418 493
<< viali >>
rect 3374 2449 3408 2483
rect 798 2247 832 2281
rect 1409 2247 1443 2281
rect 1627 2247 1661 2281
rect 2237 2247 2271 2281
rect 2548 2247 2582 2281
rect 3170 2247 3204 2281
rect 1250 1871 1284 1905
rect 847 1783 881 1817
rect 937 1783 971 1817
rect 1079 1783 1113 1817
rect 1247 1783 1281 1817
rect 1491 1783 1525 1817
rect 1581 1783 1615 1817
rect 1767 1783 1801 1817
rect 1857 1784 1891 1818
rect 2000 1783 2034 1817
rect 2353 1783 2387 1817
rect 2574 1783 2608 1817
rect 3183 1783 3217 1817
rect 3308 1471 3342 1505
rect 805 1159 839 1193
rect 973 1159 1007 1193
rect 1307 1159 1341 1193
rect 1396 1159 1430 1193
rect 1767 1159 1801 1193
rect 1857 1159 1891 1193
rect 2000 1159 2034 1193
rect 2356 1159 2390 1193
rect 2574 1159 2608 1193
rect 3184 1159 3218 1193
rect 802 1071 836 1105
rect 705 927 739 961
rect 796 695 830 729
rect 1409 695 1443 729
rect 1627 695 1661 729
rect 2237 695 2271 729
rect 2546 695 2580 729
rect 3156 695 3190 729
rect 3360 493 3394 527
<< metal1 >>
rect 2423 2528 2514 2624
rect 3299 2528 3550 2624
rect 3343 2483 3550 2528
rect 3343 2449 3374 2483
rect 3408 2449 3550 2483
rect 3343 2418 3550 2449
rect 748 2281 844 2287
rect 748 2247 798 2281
rect 832 2247 844 2281
rect 748 2241 844 2247
rect 1397 2281 1673 2287
rect 1397 2247 1409 2281
rect 1443 2247 1627 2281
rect 1661 2247 1673 2281
rect 1397 2241 1673 2247
rect 2225 2281 2594 2287
rect 2225 2247 2237 2281
rect 2271 2247 2548 2281
rect 2582 2247 2594 2281
rect 2225 2241 2594 2247
rect 3158 2281 3415 2287
rect 3158 2247 3170 2281
rect 3204 2247 3415 2281
rect 3158 2241 3415 2247
rect 565 1984 842 2080
rect 565 992 661 1984
rect 3374 1942 3415 2241
rect 1238 1905 1449 1911
rect 1238 1871 1250 1905
rect 1284 1871 1449 1905
rect 3362 1890 3368 1942
rect 3420 1890 3426 1942
rect 1238 1865 1449 1871
rect 1403 1823 1449 1865
rect 689 1817 893 1823
rect 689 1783 847 1817
rect 881 1783 893 1817
rect 689 1777 893 1783
rect 925 1817 1125 1823
rect 925 1783 937 1817
rect 971 1783 1079 1817
rect 1113 1783 1125 1817
rect 925 1777 1125 1783
rect 1235 1817 1365 1823
rect 1235 1783 1247 1817
rect 1281 1783 1365 1817
rect 1235 1777 1365 1783
rect 1403 1817 1537 1823
rect 1403 1783 1491 1817
rect 1525 1783 1537 1817
rect 1403 1777 1537 1783
rect 1569 1817 1813 1823
rect 1569 1783 1581 1817
rect 1615 1783 1767 1817
rect 1801 1783 1813 1817
rect 1569 1777 1813 1783
rect 1845 1818 2046 1824
rect 3374 1823 3415 1890
rect 1845 1784 1857 1818
rect 1891 1817 2046 1818
rect 1891 1784 2000 1817
rect 1845 1783 2000 1784
rect 2034 1783 2046 1817
rect 1845 1777 2046 1783
rect 2341 1817 2620 1823
rect 2341 1783 2353 1817
rect 2387 1783 2574 1817
rect 2608 1783 2620 1817
rect 2341 1777 2620 1783
rect 3171 1817 3415 1823
rect 3171 1783 3183 1817
rect 3217 1783 3415 1817
rect 3171 1777 3415 1783
rect 689 1199 739 1777
rect 1318 1695 1365 1777
rect 1318 1686 1417 1695
rect 1318 1634 1365 1686
rect 1417 1634 1423 1686
rect 3454 1536 3550 2418
rect 3232 1505 3550 1536
rect 3232 1471 3308 1505
rect 3342 1471 3550 1505
rect 3232 1440 3550 1471
rect 3283 1399 3335 1405
rect 1011 1269 1017 1321
rect 1069 1269 1075 1321
rect 1020 1199 1066 1269
rect 689 1193 851 1199
rect 689 1159 805 1193
rect 839 1159 851 1193
rect 689 1153 851 1159
rect 961 1193 1066 1199
rect 961 1159 973 1193
rect 1007 1159 1066 1193
rect 961 1153 1066 1159
rect 1101 1150 1107 1202
rect 1159 1199 1165 1202
rect 1159 1193 1353 1199
rect 1159 1159 1307 1193
rect 1341 1159 1353 1193
rect 1159 1153 1353 1159
rect 1384 1193 1813 1199
rect 1384 1159 1396 1193
rect 1430 1159 1767 1193
rect 1801 1159 1813 1193
rect 1384 1153 1813 1159
rect 1845 1193 2046 1199
rect 1845 1159 1857 1193
rect 1891 1159 2000 1193
rect 2034 1159 2046 1193
rect 1845 1153 2046 1159
rect 2344 1193 2620 1206
rect 3283 1199 3335 1347
rect 2344 1159 2356 1193
rect 2390 1159 2574 1193
rect 2608 1159 2620 1193
rect 2344 1153 2620 1159
rect 3172 1193 3335 1199
rect 3172 1159 3184 1193
rect 3218 1159 3335 1193
rect 3172 1153 3335 1159
rect 1159 1150 1165 1153
rect 707 1114 759 1120
rect 759 1105 848 1111
rect 759 1071 802 1105
rect 836 1071 848 1105
rect 759 1065 848 1071
rect 3283 1088 3335 1153
rect 707 1056 759 1062
rect 3283 1030 3335 1036
rect 565 961 787 992
rect 565 927 705 961
rect 739 927 790 961
rect 565 896 787 927
rect 3260 895 3317 896
rect 3283 735 3335 737
rect 758 729 848 735
rect 758 695 796 729
rect 830 695 848 729
rect 758 685 848 695
rect 1397 729 1673 735
rect 1397 695 1409 729
rect 1443 695 1627 729
rect 1661 695 1673 729
rect 1397 689 1673 695
rect 2225 729 2592 735
rect 2225 695 2237 729
rect 2271 695 2546 729
rect 2580 695 2592 729
rect 2225 689 2592 695
rect 3144 731 3335 735
rect 3144 729 3283 731
rect 3144 695 3156 729
rect 3190 695 3283 729
rect 3144 679 3283 695
rect 3283 673 3335 679
rect 3454 558 3550 1440
rect 3329 527 3550 558
rect 3329 493 3360 527
rect 3394 493 3550 527
rect 3329 448 3550 493
rect 2423 352 2514 448
rect 3314 352 3550 448
<< via1 >>
rect 3368 1890 3420 1942
rect 1365 1634 1417 1686
rect 3283 1347 3335 1399
rect 1017 1269 1069 1321
rect 1107 1150 1159 1202
rect 707 1062 759 1114
rect 3283 1036 3335 1088
rect 3283 679 3335 731
<< metal2 >>
rect 995 2009 3419 2055
rect 995 1593 1041 2009
rect 3369 1948 3419 2009
rect 3368 1942 3420 1948
rect 3368 1884 3420 1890
rect 1365 1686 1417 1695
rect 995 1544 1066 1593
rect 1020 1327 1066 1544
rect 1365 1505 1417 1634
rect 1365 1470 3335 1505
rect 3283 1399 3335 1470
rect 3277 1347 3283 1399
rect 3335 1347 3341 1399
rect 1017 1321 1069 1327
rect 1017 1263 1069 1269
rect 1107 1202 1159 1208
rect 1107 1144 1159 1150
rect 701 1062 707 1114
rect 759 1062 765 1114
rect 710 970 756 1062
rect 1109 970 1157 1144
rect 3277 1036 3283 1088
rect 3335 1036 3341 1088
rect 710 924 1157 970
rect 1109 923 1157 924
rect 3283 731 3335 1036
rect 3277 679 3283 731
rect 3335 679 3341 731
use sky130_fd_sc_hd__nand2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1043 0 1 944
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x2
timestamp 1704896540
transform 1 0 1043 0 -1 2032
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 767 0 -1 2032
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4
timestamp 1704896540
transform 1 0 1227 0 1 944
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1704896540
transform 1 0 1411 0 -1 2032
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1704896540
transform 1 0 1687 0 1 944
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1704896540
transform 1 0 1687 0 -1 2032
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1963 0 1 944
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  x9
timestamp 1704896540
transform 1 0 1963 0 -1 2032
box -38 -48 498 592
use sky130_fd_sc_hd__inv_8  x10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2423 0 -1 944
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x11
timestamp 1704896540
transform -1 0 2423 0 1 2032
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x12
timestamp 1704896540
transform -1 0 1595 0 -1 944
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x13
timestamp 1704896540
transform -1 0 1595 0 1 2032
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x14
timestamp 1704896540
transform 1 0 2422 0 1 944
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x15
timestamp 1704896540
transform 1 0 2422 0 -1 2032
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x16
timestamp 1704896540
transform 1 0 2514 0 1 2032
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x17
timestamp 1704896540
transform -1 0 3342 0 -1 944
box -38 -48 866 592
<< labels >>
flabel metal1 3415 1482 3415 1482 0 FreeSans 800 0 0 0 VDDA
port 0 nsew
flabel metal1 606 1478 606 1478 0 FreeSans 800 0 0 0 VSSA
port 1 nsew
flabel metal1 722 1184 722 1184 0 FreeSans 800 0 0 0 in
port 2 nsew
flabel metal1 767 709 767 709 0 FreeSans 800 0 0 0 clk0
port 3 nsew
flabel metal1 764 2262 764 2262 0 FreeSans 800 0 0 0 clk1
port 4 nsew
flabel metal1 1588 709 1589 709 0 FreeSans 800 0 0 0 clkb0
port 5 nsew
flabel metal1 1592 2265 1593 2265 0 FreeSans 800 0 0 0 clkb1
port 6 nsew
<< end >>
