magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 1 21 1715 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 177 47 207 177
rect 271 47 301 177
rect 375 47 405 177
rect 459 47 489 177
rect 553 47 583 177
rect 647 47 677 177
rect 751 47 781 177
rect 939 47 969 177
rect 1033 47 1063 177
rect 1127 47 1157 177
rect 1231 47 1261 177
rect 1315 47 1345 177
rect 1409 47 1439 177
rect 1503 47 1533 177
rect 1607 47 1637 177
<< scpmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 461 297 497 497
rect 555 297 591 497
rect 649 297 685 497
rect 743 297 779 497
rect 941 297 977 497
rect 1035 297 1071 497
rect 1129 297 1165 497
rect 1223 297 1259 497
rect 1317 297 1353 497
rect 1411 297 1447 497
rect 1505 297 1541 497
rect 1599 297 1635 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 177 177
rect 113 129 133 163
rect 167 129 177 163
rect 113 95 177 129
rect 113 61 133 95
rect 167 61 177 95
rect 113 47 177 61
rect 207 95 271 177
rect 207 61 227 95
rect 261 61 271 95
rect 207 47 271 61
rect 301 163 375 177
rect 301 129 321 163
rect 355 129 375 163
rect 301 95 375 129
rect 301 61 321 95
rect 355 61 375 95
rect 301 47 375 61
rect 405 95 459 177
rect 405 61 415 95
rect 449 61 459 95
rect 405 47 459 61
rect 489 163 553 177
rect 489 129 509 163
rect 543 129 553 163
rect 489 95 553 129
rect 489 61 509 95
rect 543 61 553 95
rect 489 47 553 61
rect 583 95 647 177
rect 583 61 603 95
rect 637 61 647 95
rect 583 47 647 61
rect 677 163 751 177
rect 677 129 697 163
rect 731 129 751 163
rect 677 95 751 129
rect 677 61 697 95
rect 731 61 751 95
rect 677 47 751 61
rect 781 95 939 177
rect 781 61 791 95
rect 825 61 895 95
rect 929 61 939 95
rect 781 47 939 61
rect 969 163 1033 177
rect 969 129 989 163
rect 1023 129 1033 163
rect 969 95 1033 129
rect 969 61 989 95
rect 1023 61 1033 95
rect 969 47 1033 61
rect 1063 95 1127 177
rect 1063 61 1083 95
rect 1117 61 1127 95
rect 1063 47 1127 61
rect 1157 163 1231 177
rect 1157 129 1177 163
rect 1211 129 1231 163
rect 1157 95 1231 129
rect 1157 61 1177 95
rect 1211 61 1231 95
rect 1157 47 1231 61
rect 1261 95 1315 177
rect 1261 61 1271 95
rect 1305 61 1315 95
rect 1261 47 1315 61
rect 1345 163 1409 177
rect 1345 129 1365 163
rect 1399 129 1409 163
rect 1345 95 1409 129
rect 1345 61 1365 95
rect 1399 61 1409 95
rect 1345 47 1409 61
rect 1439 95 1503 177
rect 1439 61 1459 95
rect 1493 61 1503 95
rect 1439 47 1503 61
rect 1533 163 1607 177
rect 1533 129 1553 163
rect 1587 129 1607 163
rect 1533 95 1607 129
rect 1533 61 1553 95
rect 1587 61 1607 95
rect 1533 47 1607 61
rect 1637 95 1689 177
rect 1637 61 1647 95
rect 1681 61 1689 95
rect 1637 47 1689 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 297 179 375
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 477 367 497
rect 309 443 321 477
rect 355 443 367 477
rect 309 409 367 443
rect 309 375 321 409
rect 355 375 367 409
rect 309 297 367 375
rect 403 477 461 497
rect 403 443 415 477
rect 449 443 461 477
rect 403 409 461 443
rect 403 375 415 409
rect 449 375 461 409
rect 403 341 461 375
rect 403 307 415 341
rect 449 307 461 341
rect 403 297 461 307
rect 497 409 555 497
rect 497 375 509 409
rect 543 375 555 409
rect 497 341 555 375
rect 497 307 509 341
rect 543 307 555 341
rect 497 297 555 307
rect 591 477 649 497
rect 591 443 603 477
rect 637 443 649 477
rect 591 409 649 443
rect 591 375 603 409
rect 637 375 649 409
rect 591 297 649 375
rect 685 409 743 497
rect 685 375 697 409
rect 731 375 743 409
rect 685 341 743 375
rect 685 307 697 341
rect 731 307 743 341
rect 685 297 743 307
rect 779 477 833 497
rect 779 443 791 477
rect 825 443 833 477
rect 779 409 833 443
rect 779 375 791 409
rect 825 375 833 409
rect 779 297 833 375
rect 887 477 941 497
rect 887 443 895 477
rect 929 443 941 477
rect 887 409 941 443
rect 887 375 895 409
rect 929 375 941 409
rect 887 297 941 375
rect 977 409 1035 497
rect 977 375 989 409
rect 1023 375 1035 409
rect 977 341 1035 375
rect 977 307 989 341
rect 1023 307 1035 341
rect 977 297 1035 307
rect 1071 477 1129 497
rect 1071 443 1083 477
rect 1117 443 1129 477
rect 1071 409 1129 443
rect 1071 375 1083 409
rect 1117 375 1129 409
rect 1071 297 1129 375
rect 1165 409 1223 497
rect 1165 375 1177 409
rect 1211 375 1223 409
rect 1165 341 1223 375
rect 1165 307 1177 341
rect 1211 307 1223 341
rect 1165 297 1223 307
rect 1259 477 1317 497
rect 1259 443 1271 477
rect 1305 443 1317 477
rect 1259 409 1317 443
rect 1259 375 1271 409
rect 1305 375 1317 409
rect 1259 297 1317 375
rect 1353 409 1411 497
rect 1353 375 1365 409
rect 1399 375 1411 409
rect 1353 341 1411 375
rect 1353 307 1365 341
rect 1399 307 1411 341
rect 1353 297 1411 307
rect 1447 477 1505 497
rect 1447 443 1459 477
rect 1493 443 1505 477
rect 1447 409 1505 443
rect 1447 375 1459 409
rect 1493 375 1505 409
rect 1447 297 1505 375
rect 1541 409 1599 497
rect 1541 375 1553 409
rect 1587 375 1599 409
rect 1541 341 1599 375
rect 1541 307 1553 341
rect 1587 307 1599 341
rect 1541 297 1599 307
rect 1635 477 1689 497
rect 1635 443 1647 477
rect 1681 443 1689 477
rect 1635 409 1689 443
rect 1635 375 1647 409
rect 1681 375 1689 409
rect 1635 297 1689 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 415 61 449 95
rect 509 129 543 163
rect 509 61 543 95
rect 603 61 637 95
rect 697 129 731 163
rect 697 61 731 95
rect 791 61 825 95
rect 895 61 929 95
rect 989 129 1023 163
rect 989 61 1023 95
rect 1083 61 1117 95
rect 1177 129 1211 163
rect 1177 61 1211 95
rect 1271 61 1305 95
rect 1365 129 1399 163
rect 1365 61 1399 95
rect 1459 61 1493 95
rect 1553 129 1587 163
rect 1553 61 1587 95
rect 1647 61 1681 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 443 167 477
rect 133 375 167 409
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 443 355 477
rect 321 375 355 409
rect 415 443 449 477
rect 415 375 449 409
rect 415 307 449 341
rect 509 375 543 409
rect 509 307 543 341
rect 603 443 637 477
rect 603 375 637 409
rect 697 375 731 409
rect 697 307 731 341
rect 791 443 825 477
rect 791 375 825 409
rect 895 443 929 477
rect 895 375 929 409
rect 989 375 1023 409
rect 989 307 1023 341
rect 1083 443 1117 477
rect 1083 375 1117 409
rect 1177 375 1211 409
rect 1177 307 1211 341
rect 1271 443 1305 477
rect 1271 375 1305 409
rect 1365 375 1399 409
rect 1365 307 1399 341
rect 1459 443 1493 477
rect 1459 375 1493 409
rect 1553 375 1587 409
rect 1553 307 1587 341
rect 1647 443 1681 477
rect 1647 375 1681 409
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 461 497 497 523
rect 555 497 591 523
rect 649 497 685 523
rect 743 497 779 523
rect 941 497 977 523
rect 1035 497 1071 523
rect 1129 497 1165 523
rect 1223 497 1259 523
rect 1317 497 1353 523
rect 1411 497 1447 523
rect 1505 497 1541 523
rect 1599 497 1635 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 461 282 497 297
rect 555 282 591 297
rect 649 282 685 297
rect 743 282 779 297
rect 941 282 977 297
rect 1035 282 1071 297
rect 1129 282 1165 297
rect 1223 282 1259 297
rect 1317 282 1353 297
rect 1411 282 1447 297
rect 1505 282 1541 297
rect 1599 282 1635 297
rect 83 265 123 282
rect 177 265 217 282
rect 271 265 311 282
rect 365 265 405 282
rect 83 249 405 265
rect 83 215 99 249
rect 133 215 177 249
rect 211 215 255 249
rect 289 215 333 249
rect 367 215 405 249
rect 83 199 405 215
rect 83 177 113 199
rect 177 177 207 199
rect 271 177 301 199
rect 375 177 405 199
rect 459 265 499 282
rect 553 265 593 282
rect 647 265 687 282
rect 741 265 781 282
rect 459 249 781 265
rect 459 215 475 249
rect 509 215 553 249
rect 587 215 631 249
rect 665 215 709 249
rect 743 215 781 249
rect 459 199 781 215
rect 459 177 489 199
rect 553 177 583 199
rect 647 177 677 199
rect 751 177 781 199
rect 939 265 979 282
rect 1033 265 1073 282
rect 1127 265 1167 282
rect 1221 265 1261 282
rect 939 249 1261 265
rect 939 215 955 249
rect 989 215 1033 249
rect 1067 215 1111 249
rect 1145 215 1189 249
rect 1223 215 1261 249
rect 939 199 1261 215
rect 939 177 969 199
rect 1033 177 1063 199
rect 1127 177 1157 199
rect 1231 177 1261 199
rect 1315 265 1355 282
rect 1409 265 1449 282
rect 1503 265 1543 282
rect 1597 265 1637 282
rect 1315 249 1637 265
rect 1315 215 1325 249
rect 1359 215 1403 249
rect 1437 215 1481 249
rect 1515 215 1559 249
rect 1593 215 1637 249
rect 1315 199 1637 215
rect 1315 177 1345 199
rect 1409 177 1439 199
rect 1503 177 1533 199
rect 1607 177 1637 199
rect 83 21 113 47
rect 177 21 207 47
rect 271 21 301 47
rect 375 21 405 47
rect 459 21 489 47
rect 553 21 583 47
rect 647 21 677 47
rect 751 21 781 47
rect 939 21 969 47
rect 1033 21 1063 47
rect 1127 21 1157 47
rect 1231 21 1261 47
rect 1315 21 1345 47
rect 1409 21 1439 47
rect 1503 21 1533 47
rect 1607 21 1637 47
<< polycont >>
rect 99 215 133 249
rect 177 215 211 249
rect 255 215 289 249
rect 333 215 367 249
rect 475 215 509 249
rect 553 215 587 249
rect 631 215 665 249
rect 709 215 743 249
rect 955 215 989 249
rect 1033 215 1067 249
rect 1111 215 1145 249
rect 1189 215 1223 249
rect 1325 215 1359 249
rect 1403 215 1437 249
rect 1481 215 1515 249
rect 1559 215 1593 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 18 477 81 493
rect 18 443 39 477
rect 73 443 81 477
rect 18 409 81 443
rect 18 375 39 409
rect 73 375 81 409
rect 18 341 81 375
rect 125 477 175 527
rect 125 443 133 477
rect 167 443 175 477
rect 125 409 175 443
rect 125 375 133 409
rect 167 375 175 409
rect 125 359 175 375
rect 219 477 269 493
rect 219 443 227 477
rect 261 443 269 477
rect 219 409 269 443
rect 219 375 227 409
rect 261 375 269 409
rect 18 307 39 341
rect 73 325 81 341
rect 219 341 269 375
rect 313 477 363 527
rect 313 443 321 477
rect 355 443 363 477
rect 313 409 363 443
rect 313 375 321 409
rect 355 375 363 409
rect 313 359 363 375
rect 407 477 844 493
rect 407 443 415 477
rect 449 459 603 477
rect 449 443 457 459
rect 407 409 457 443
rect 595 443 603 459
rect 637 459 791 477
rect 637 443 645 459
rect 407 375 415 409
rect 449 375 457 409
rect 219 325 227 341
rect 73 307 227 325
rect 261 325 269 341
rect 407 341 457 375
rect 407 325 415 341
rect 261 307 415 325
rect 449 307 457 341
rect 18 291 457 307
rect 501 409 551 425
rect 501 375 509 409
rect 543 375 551 409
rect 501 341 551 375
rect 595 409 645 443
rect 783 443 791 459
rect 825 443 844 477
rect 595 375 603 409
rect 637 375 645 409
rect 595 359 645 375
rect 689 409 739 425
rect 689 375 697 409
rect 731 375 739 409
rect 501 307 509 341
rect 543 325 551 341
rect 689 341 739 375
rect 783 409 844 443
rect 783 375 791 409
rect 825 375 844 409
rect 783 359 844 375
rect 881 477 1689 493
rect 881 443 895 477
rect 929 459 1083 477
rect 929 443 937 459
rect 881 409 937 443
rect 1075 443 1083 459
rect 1117 459 1271 477
rect 1117 443 1125 459
rect 881 375 895 409
rect 929 375 937 409
rect 881 359 937 375
rect 981 409 1031 425
rect 981 375 989 409
rect 1023 375 1031 409
rect 689 325 697 341
rect 543 307 697 325
rect 731 325 739 341
rect 981 341 1031 375
rect 1075 409 1125 443
rect 1263 443 1271 459
rect 1305 459 1459 477
rect 1305 443 1313 459
rect 1075 375 1083 409
rect 1117 375 1125 409
rect 1075 359 1125 375
rect 1169 409 1219 425
rect 1169 375 1177 409
rect 1211 375 1219 409
rect 981 325 989 341
rect 731 307 989 325
rect 1023 325 1031 341
rect 1169 341 1219 375
rect 1263 409 1313 443
rect 1451 443 1459 459
rect 1493 459 1647 477
rect 1493 443 1501 459
rect 1263 375 1271 409
rect 1305 375 1313 409
rect 1263 359 1313 375
rect 1357 409 1407 425
rect 1357 375 1365 409
rect 1399 375 1407 409
rect 1169 325 1177 341
rect 1023 307 1177 325
rect 1211 307 1219 341
rect 501 291 1219 307
rect 1357 341 1407 375
rect 1451 409 1501 443
rect 1639 443 1647 459
rect 1681 443 1689 477
rect 1451 375 1459 409
rect 1493 375 1501 409
rect 1451 359 1501 375
rect 1545 409 1595 425
rect 1545 375 1553 409
rect 1587 375 1595 409
rect 1357 307 1365 341
rect 1399 325 1407 341
rect 1545 341 1595 375
rect 1639 409 1689 443
rect 1639 375 1647 409
rect 1681 375 1689 409
rect 1639 359 1689 375
rect 1545 325 1553 341
rect 1399 307 1553 325
rect 1587 325 1595 341
rect 1587 307 1726 325
rect 1357 291 1726 307
rect 36 249 405 257
rect 36 215 99 249
rect 133 215 177 249
rect 211 215 255 249
rect 289 215 333 249
rect 367 215 405 249
rect 459 249 894 257
rect 459 215 475 249
rect 509 215 553 249
rect 587 215 631 249
rect 665 215 709 249
rect 743 215 894 249
rect 939 249 1261 257
rect 939 215 955 249
rect 989 215 1033 249
rect 1067 215 1111 249
rect 1145 215 1189 249
rect 1223 215 1261 249
rect 1295 249 1609 257
rect 1295 215 1325 249
rect 1359 215 1403 249
rect 1437 215 1481 249
rect 1515 215 1559 249
rect 1593 215 1609 249
rect 1672 181 1726 291
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 1726 181
rect 107 129 133 163
rect 167 145 321 163
rect 167 129 183 145
rect 107 95 183 129
rect 295 129 321 145
rect 355 145 509 163
rect 355 129 371 145
rect 107 61 133 95
rect 167 61 183 95
rect 107 51 183 61
rect 227 95 261 111
rect 227 17 261 61
rect 295 95 371 129
rect 483 129 509 145
rect 543 145 697 163
rect 543 129 559 145
rect 295 61 321 95
rect 355 61 371 95
rect 295 51 371 61
rect 415 95 449 111
rect 415 17 449 61
rect 483 95 559 129
rect 671 129 697 145
rect 731 145 989 163
rect 731 129 747 145
rect 483 61 509 95
rect 543 61 559 95
rect 483 51 559 61
rect 603 95 637 111
rect 603 17 637 61
rect 671 95 747 129
rect 963 129 989 145
rect 1023 145 1177 163
rect 1023 129 1039 145
rect 671 61 697 95
rect 731 61 747 95
rect 671 51 747 61
rect 791 95 929 111
rect 825 61 895 95
rect 791 17 929 61
rect 963 95 1039 129
rect 1151 129 1177 145
rect 1211 145 1365 163
rect 1211 129 1227 145
rect 963 61 989 95
rect 1023 61 1039 95
rect 963 51 1039 61
rect 1083 95 1117 111
rect 1083 17 1117 61
rect 1151 95 1227 129
rect 1339 129 1365 145
rect 1399 145 1553 163
rect 1399 129 1415 145
rect 1151 61 1177 95
rect 1211 61 1227 95
rect 1151 51 1227 61
rect 1271 95 1305 111
rect 1271 17 1305 61
rect 1339 95 1415 129
rect 1527 129 1553 145
rect 1587 145 1726 163
rect 1587 129 1603 145
rect 1339 61 1365 95
rect 1399 61 1415 95
rect 1339 51 1415 61
rect 1459 95 1493 111
rect 1459 17 1493 61
rect 1527 95 1603 129
rect 1527 61 1553 95
rect 1587 61 1603 95
rect 1527 51 1603 61
rect 1647 95 1681 111
rect 1647 17 1681 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel locali s 36 215 405 257 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 1040 221 1074 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 1672 181 1726 291 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 1458 221 1492 255 0 FreeSans 400 0 0 0 D
port 4 nsew signal input
flabel locali s 846 221 880 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 744 221 778 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 642 221 676 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4_4
rlabel locali s 1545 325 1595 425 1 Y
port 9 nsew signal output
rlabel locali s 1527 51 1603 145 1 Y
port 9 nsew signal output
rlabel locali s 1357 325 1407 425 1 Y
port 9 nsew signal output
rlabel locali s 1357 291 1726 325 1 Y
port 9 nsew signal output
rlabel locali s 1339 51 1415 145 1 Y
port 9 nsew signal output
rlabel locali s 1151 51 1227 145 1 Y
port 9 nsew signal output
rlabel locali s 963 51 1039 145 1 Y
port 9 nsew signal output
rlabel locali s 671 51 747 145 1 Y
port 9 nsew signal output
rlabel locali s 483 51 559 145 1 Y
port 9 nsew signal output
rlabel locali s 295 51 371 145 1 Y
port 9 nsew signal output
rlabel locali s 107 145 1726 181 1 Y
port 9 nsew signal output
rlabel locali s 107 51 183 145 1 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_END 1789634
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1776516
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
