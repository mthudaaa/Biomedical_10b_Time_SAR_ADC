magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 157 197 203
rect 1 21 881 157
rect 84 -17 128 21
<< scnmos >>
rect 79 47 109 177
rect 215 47 245 131
rect 317 47 347 131
rect 469 47 499 131
rect 657 47 687 131
rect 773 47 803 131
<< scpmoshvt >>
rect 81 297 117 497
rect 207 374 243 458
rect 326 374 362 458
rect 577 374 613 458
rect 659 374 695 458
rect 765 374 801 458
<< ndiff >>
rect 27 112 79 177
rect 27 78 35 112
rect 69 78 79 112
rect 27 47 79 78
rect 109 131 171 177
rect 109 93 215 131
rect 109 59 129 93
rect 163 59 215 93
rect 109 47 215 59
rect 245 47 317 131
rect 347 108 469 131
rect 347 74 357 108
rect 391 74 469 108
rect 347 47 469 74
rect 499 47 657 131
rect 687 108 773 131
rect 687 74 719 108
rect 753 74 773 108
rect 687 47 773 74
rect 803 108 855 131
rect 803 74 813 108
rect 847 74 855 108
rect 803 47 855 74
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 171 497
rect 117 451 129 485
rect 163 458 171 485
rect 163 451 207 458
rect 117 417 207 451
rect 117 383 129 417
rect 163 383 207 417
rect 117 374 207 383
rect 243 374 326 458
rect 362 425 577 458
rect 362 391 385 425
rect 419 391 490 425
rect 524 391 577 425
rect 362 374 577 391
rect 613 374 659 458
rect 695 425 765 458
rect 695 391 717 425
rect 751 391 765 425
rect 695 374 765 391
rect 801 425 859 458
rect 801 391 813 425
rect 847 391 859 425
rect 801 374 859 391
rect 117 349 171 374
rect 117 315 129 349
rect 163 315 171 349
rect 117 297 171 315
<< ndiffc >>
rect 35 78 69 112
rect 129 59 163 93
rect 357 74 391 108
rect 719 74 753 108
rect 813 74 847 108
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 385 391 419 425
rect 490 391 524 425
rect 717 391 751 425
rect 813 391 847 425
rect 129 315 163 349
<< poly >>
rect 81 497 117 523
rect 207 458 243 484
rect 326 458 362 484
rect 577 458 613 484
rect 659 458 695 484
rect 765 458 801 484
rect 207 359 243 374
rect 326 359 362 374
rect 577 359 613 374
rect 659 359 695 374
rect 765 359 801 374
rect 81 282 117 297
rect 79 265 119 282
rect 205 265 245 359
rect 324 329 509 359
rect 575 342 615 359
rect 79 249 147 265
rect 79 215 103 249
rect 137 215 147 249
rect 79 199 147 215
rect 189 249 245 265
rect 189 215 199 249
rect 233 215 245 249
rect 469 229 509 329
rect 561 326 615 342
rect 561 292 571 326
rect 605 292 615 326
rect 561 276 615 292
rect 189 199 245 215
rect 79 177 109 199
rect 215 131 245 199
rect 317 213 400 229
rect 317 179 356 213
rect 390 179 400 213
rect 317 163 400 179
rect 469 213 533 229
rect 469 179 479 213
rect 513 179 533 213
rect 469 163 533 179
rect 657 223 697 359
rect 763 342 803 359
rect 739 326 803 342
rect 739 292 749 326
rect 783 292 803 326
rect 739 276 803 292
rect 657 213 723 223
rect 657 179 673 213
rect 707 179 723 213
rect 657 169 723 179
rect 317 131 347 163
rect 469 131 499 163
rect 657 131 687 169
rect 773 131 803 276
rect 79 21 109 47
rect 215 21 245 47
rect 317 21 347 47
rect 469 21 499 47
rect 657 21 687 47
rect 773 21 803 47
<< polycont >>
rect 103 215 137 249
rect 199 215 233 249
rect 571 292 605 326
rect 356 179 390 213
rect 479 179 513 213
rect 749 292 783 326
rect 673 179 707 213
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 485 85 493
rect 18 451 35 485
rect 69 451 85 485
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 18 349 85 383
rect 18 315 35 349
rect 69 315 85 349
rect 18 299 85 315
rect 129 485 163 527
rect 129 417 163 451
rect 129 349 163 383
rect 129 299 163 315
rect 214 459 683 493
rect 18 112 69 299
rect 214 265 254 459
rect 103 249 137 265
rect 103 165 137 215
rect 199 249 254 265
rect 233 215 254 249
rect 199 199 254 215
rect 288 391 385 425
rect 419 391 490 425
rect 524 391 550 425
rect 288 165 322 391
rect 103 131 322 165
rect 356 326 615 357
rect 356 323 571 326
rect 356 213 390 323
rect 605 292 615 326
rect 356 163 390 179
rect 458 213 523 283
rect 458 179 479 213
rect 513 179 523 213
rect 18 78 35 112
rect 287 124 322 131
rect 287 108 391 124
rect 18 51 69 78
rect 103 93 179 97
rect 103 59 129 93
rect 163 59 179 93
rect 103 17 179 59
rect 287 74 357 108
rect 287 51 391 74
rect 458 51 523 179
rect 571 51 615 292
rect 649 326 683 459
rect 717 425 751 527
rect 717 375 751 391
rect 808 425 900 457
rect 808 391 813 425
rect 847 391 900 425
rect 808 375 900 391
rect 649 292 749 326
rect 783 292 809 326
rect 649 288 809 292
rect 843 213 900 375
rect 657 179 673 213
rect 707 179 900 213
rect 650 108 753 124
rect 650 74 719 108
rect 650 17 753 74
rect 807 108 856 179
rect 807 74 813 108
rect 847 74 856 108
rect 807 58 856 74
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
flabel locali s 672 289 706 323 0 FreeSans 250 0 0 0 S
port 3 nsew signal input
flabel locali s 579 153 613 187 0 FreeSans 250 0 0 0 A1
port 2 nsew signal input
flabel locali s 577 221 611 255 0 FreeSans 250 0 0 0 A1
port 2 nsew signal input
flabel locali s 458 51 523 283 0 FreeSans 250 0 0 0 A0
port 1 nsew signal input
flabel locali s 30 85 64 119 0 FreeSans 250 0 0 0 X
port 8 nsew signal output
flabel locali s 30 357 64 391 0 FreeSans 250 0 0 0 X
port 8 nsew signal output
flabel locali s 30 425 64 459 0 FreeSans 250 0 0 0 X
port 8 nsew signal output
flabel locali s 761 289 795 323 0 FreeSans 250 0 0 0 S
port 3 nsew signal input
flabel nwell s 74 527 108 561 0 FreeSans 250 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 84 -17 128 17 0 FreeSans 250 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 mux2_1
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 1417444
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1410552
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
