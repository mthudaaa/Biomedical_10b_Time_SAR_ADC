magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 723 203
rect 30 -17 64 21
<< scnmos >>
rect 80 47 110 177
rect 196 47 226 177
rect 374 47 404 177
rect 502 47 532 177
rect 605 47 635 177
<< scpmoshvt >>
rect 82 297 118 497
rect 188 297 224 497
rect 408 297 444 497
rect 504 297 540 497
rect 607 297 643 497
<< ndiff >>
rect 27 93 80 177
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 101 196 177
rect 110 67 131 101
rect 165 67 196 101
rect 110 47 196 67
rect 226 89 374 177
rect 226 55 281 89
rect 315 55 374 89
rect 226 47 374 55
rect 404 101 502 177
rect 404 67 414 101
rect 448 67 502 101
rect 404 47 502 67
rect 532 47 605 177
rect 635 93 697 177
rect 635 59 655 93
rect 689 59 697 93
rect 635 47 697 59
<< pdiff >>
rect 27 485 82 497
rect 27 451 35 485
rect 69 451 82 485
rect 27 386 82 451
rect 27 352 35 386
rect 69 352 82 386
rect 27 297 82 352
rect 118 477 188 497
rect 118 443 131 477
rect 165 443 188 477
rect 118 382 188 443
rect 118 348 131 382
rect 165 348 188 382
rect 118 297 188 348
rect 224 485 289 497
rect 224 451 237 485
rect 271 451 289 485
rect 224 297 289 451
rect 343 477 408 497
rect 343 443 351 477
rect 385 443 408 477
rect 343 393 408 443
rect 343 359 351 393
rect 385 359 408 393
rect 343 297 408 359
rect 444 477 504 497
rect 444 443 457 477
rect 491 443 504 477
rect 444 387 504 443
rect 444 353 457 387
rect 491 353 504 387
rect 444 297 504 353
rect 540 485 607 497
rect 540 451 557 485
rect 591 451 607 485
rect 540 297 607 451
rect 643 477 697 497
rect 643 443 655 477
rect 689 443 697 477
rect 643 387 697 443
rect 643 353 655 387
rect 689 353 697 387
rect 643 297 697 353
<< ndiffc >>
rect 35 59 69 93
rect 131 67 165 101
rect 281 55 315 89
rect 414 67 448 101
rect 655 59 689 93
<< pdiffc >>
rect 35 451 69 485
rect 35 352 69 386
rect 131 443 165 477
rect 131 348 165 382
rect 237 451 271 485
rect 351 443 385 477
rect 351 359 385 393
rect 457 443 491 477
rect 457 353 491 387
rect 557 451 591 485
rect 655 443 689 477
rect 655 353 689 387
<< poly >>
rect 82 497 118 523
rect 188 497 224 523
rect 408 497 444 523
rect 504 497 540 523
rect 607 497 643 523
rect 82 282 118 297
rect 188 282 224 297
rect 408 282 444 297
rect 504 282 540 297
rect 607 282 643 297
rect 80 229 120 282
rect 186 265 226 282
rect 406 265 446 282
rect 186 249 243 265
rect 186 229 199 249
rect 80 215 199 229
rect 233 215 243 249
rect 80 199 243 215
rect 374 249 446 265
rect 374 215 394 249
rect 428 215 446 249
rect 374 199 446 215
rect 502 265 542 282
rect 605 265 645 282
rect 502 249 556 265
rect 502 215 512 249
rect 546 215 556 249
rect 502 199 556 215
rect 605 249 676 265
rect 605 215 632 249
rect 666 215 676 249
rect 605 199 676 215
rect 80 177 110 199
rect 196 177 226 199
rect 374 177 404 199
rect 502 177 532 199
rect 605 177 635 199
rect 80 21 110 47
rect 196 21 226 47
rect 374 21 404 47
rect 502 21 532 47
rect 605 21 635 47
<< polycont >>
rect 199 215 233 249
rect 394 215 428 249
rect 512 215 546 249
rect 632 215 666 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 19 485 75 527
rect 19 451 35 485
rect 69 451 75 485
rect 19 386 75 451
rect 19 352 35 386
rect 69 352 75 386
rect 19 333 75 352
rect 109 477 165 493
rect 109 443 131 477
rect 211 485 297 527
rect 211 451 237 485
rect 271 451 297 485
rect 211 444 297 451
rect 335 477 408 493
rect 109 382 165 443
rect 335 443 351 477
rect 385 443 408 477
rect 335 393 408 443
rect 335 384 351 393
rect 109 348 131 382
rect 35 93 69 111
rect 35 17 69 59
rect 109 101 165 348
rect 199 359 351 384
rect 385 359 408 393
rect 199 338 408 359
rect 452 477 497 493
rect 452 443 457 477
rect 491 443 497 477
rect 452 387 497 443
rect 541 485 607 527
rect 541 451 557 485
rect 591 451 607 485
rect 541 425 607 451
rect 651 477 695 493
rect 651 443 655 477
rect 689 443 695 477
rect 651 387 695 443
rect 452 353 457 387
rect 491 353 655 387
rect 689 353 695 387
rect 199 249 286 338
rect 452 334 695 353
rect 233 215 286 249
rect 199 165 286 215
rect 373 249 448 282
rect 373 215 394 249
rect 428 215 448 249
rect 373 199 448 215
rect 482 249 546 265
rect 482 215 512 249
rect 199 131 448 165
rect 109 67 131 101
rect 410 101 448 131
rect 109 51 165 67
rect 255 55 281 89
rect 315 55 331 89
rect 255 17 331 55
rect 410 67 414 101
rect 482 73 546 215
rect 632 249 707 265
rect 666 215 707 249
rect 632 150 707 215
rect 631 93 707 113
rect 410 51 448 67
rect 631 59 655 93
rect 689 59 707 93
rect 631 17 707 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 117 425 151 459 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 396 221 430 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 493 153 527 187 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 662 221 696 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 493 85 527 119 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21o_2
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 202550
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 196788
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
