magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1470 203
rect 29 -17 63 21
<< scnmos >>
rect 120 47 150 177
rect 226 47 256 177
rect 322 47 352 177
rect 418 47 448 177
rect 514 47 544 177
rect 694 47 724 177
rect 778 47 808 177
rect 880 47 910 177
rect 976 47 1006 177
rect 1076 47 1106 177
rect 1160 47 1190 177
rect 1264 47 1294 177
rect 1360 47 1390 177
<< scpmoshvt >>
rect 82 297 118 497
rect 292 297 328 497
rect 388 297 424 497
rect 484 297 520 497
rect 580 297 616 497
rect 682 297 718 497
rect 780 297 816 497
rect 876 297 912 497
rect 972 297 1008 497
rect 1068 297 1104 497
rect 1162 297 1198 497
rect 1256 297 1292 497
rect 1350 297 1386 497
<< ndiff >>
rect 27 157 120 177
rect 27 123 39 157
rect 73 123 120 157
rect 27 89 120 123
rect 27 55 39 89
rect 73 55 120 89
rect 27 47 120 55
rect 150 89 226 177
rect 150 55 173 89
rect 207 55 226 89
rect 150 47 226 55
rect 256 124 322 177
rect 256 90 277 124
rect 311 90 322 124
rect 256 47 322 90
rect 352 89 418 177
rect 352 55 373 89
rect 407 55 418 89
rect 352 47 418 55
rect 448 169 514 177
rect 448 135 469 169
rect 503 135 514 169
rect 448 101 514 135
rect 448 67 469 101
rect 503 67 514 101
rect 448 47 514 67
rect 544 89 694 177
rect 544 55 565 89
rect 599 55 643 89
rect 677 55 694 89
rect 544 47 694 55
rect 724 101 778 177
rect 724 67 734 101
rect 768 67 778 101
rect 724 47 778 67
rect 808 169 880 177
rect 808 135 835 169
rect 869 135 880 169
rect 808 47 880 135
rect 910 101 976 177
rect 910 67 931 101
rect 965 67 976 101
rect 910 47 976 67
rect 1006 169 1076 177
rect 1006 135 1027 169
rect 1061 135 1076 169
rect 1006 47 1076 135
rect 1106 89 1160 177
rect 1106 55 1116 89
rect 1150 55 1160 89
rect 1106 47 1160 55
rect 1190 97 1264 177
rect 1190 63 1219 97
rect 1253 63 1264 97
rect 1190 47 1264 63
rect 1294 164 1360 177
rect 1294 130 1315 164
rect 1349 130 1360 164
rect 1294 96 1360 130
rect 1294 62 1315 96
rect 1349 62 1360 96
rect 1294 47 1360 62
rect 1390 161 1444 177
rect 1390 127 1400 161
rect 1434 127 1444 161
rect 1390 93 1444 127
rect 1390 59 1400 93
rect 1434 59 1444 93
rect 1390 47 1444 59
<< pdiff >>
rect 27 485 82 497
rect 27 451 35 485
rect 69 451 82 485
rect 27 417 82 451
rect 27 383 35 417
rect 69 383 82 417
rect 27 297 82 383
rect 118 485 173 497
rect 118 451 131 485
rect 165 451 173 485
rect 118 297 173 451
rect 227 477 292 497
rect 227 443 236 477
rect 270 443 292 477
rect 227 409 292 443
rect 227 375 236 409
rect 270 375 292 409
rect 227 297 292 375
rect 328 387 388 497
rect 328 353 341 387
rect 375 353 388 387
rect 328 297 388 353
rect 424 489 484 497
rect 424 455 437 489
rect 471 455 484 489
rect 424 297 484 455
rect 520 395 580 497
rect 520 361 533 395
rect 567 361 580 395
rect 520 297 580 361
rect 616 477 682 497
rect 616 443 635 477
rect 669 443 682 477
rect 616 297 682 443
rect 718 489 780 497
rect 718 455 733 489
rect 767 455 780 489
rect 718 297 780 455
rect 816 415 876 497
rect 816 381 829 415
rect 863 381 876 415
rect 816 297 876 381
rect 912 489 972 497
rect 912 455 925 489
rect 959 455 972 489
rect 912 297 972 455
rect 1008 477 1068 497
rect 1008 443 1021 477
rect 1055 443 1068 477
rect 1008 409 1068 443
rect 1008 375 1021 409
rect 1055 375 1068 409
rect 1008 297 1068 375
rect 1104 489 1162 497
rect 1104 455 1116 489
rect 1150 455 1162 489
rect 1104 297 1162 455
rect 1198 477 1256 497
rect 1198 443 1210 477
rect 1244 443 1256 477
rect 1198 297 1256 443
rect 1292 489 1350 497
rect 1292 455 1304 489
rect 1338 455 1350 489
rect 1292 297 1350 455
rect 1386 477 1442 497
rect 1386 443 1398 477
rect 1432 443 1442 477
rect 1386 409 1442 443
rect 1386 375 1398 409
rect 1432 375 1442 409
rect 1386 297 1442 375
<< ndiffc >>
rect 39 123 73 157
rect 39 55 73 89
rect 173 55 207 89
rect 277 90 311 124
rect 373 55 407 89
rect 469 135 503 169
rect 469 67 503 101
rect 565 55 599 89
rect 643 55 677 89
rect 734 67 768 101
rect 835 135 869 169
rect 931 67 965 101
rect 1027 135 1061 169
rect 1116 55 1150 89
rect 1219 63 1253 97
rect 1315 130 1349 164
rect 1315 62 1349 96
rect 1400 127 1434 161
rect 1400 59 1434 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 131 451 165 485
rect 236 443 270 477
rect 236 375 270 409
rect 341 353 375 387
rect 437 455 471 489
rect 533 361 567 395
rect 635 443 669 477
rect 733 455 767 489
rect 829 381 863 415
rect 925 455 959 489
rect 1021 443 1055 477
rect 1021 375 1055 409
rect 1116 455 1150 489
rect 1210 443 1244 477
rect 1304 455 1338 489
rect 1398 443 1432 477
rect 1398 375 1432 409
<< poly >>
rect 82 497 118 523
rect 292 497 328 523
rect 388 497 424 523
rect 484 497 520 523
rect 580 497 616 523
rect 682 497 718 523
rect 780 497 816 523
rect 876 497 912 523
rect 972 497 1008 523
rect 1068 497 1104 523
rect 1162 497 1198 523
rect 1256 497 1292 523
rect 1350 497 1386 523
rect 82 282 118 297
rect 292 282 328 297
rect 388 282 424 297
rect 484 282 520 297
rect 580 282 616 297
rect 682 282 718 297
rect 780 282 816 297
rect 876 282 912 297
rect 972 282 1008 297
rect 1068 282 1104 297
rect 1162 282 1198 297
rect 1256 282 1292 297
rect 1350 282 1386 297
rect 80 265 120 282
rect 290 265 330 282
rect 386 265 426 282
rect 482 265 522 282
rect 578 265 618 282
rect 680 265 720 282
rect 80 249 150 265
rect 80 215 90 249
rect 124 215 150 249
rect 80 199 150 215
rect 120 177 150 199
rect 226 249 618 265
rect 226 215 292 249
rect 326 215 370 249
rect 404 215 448 249
rect 482 215 618 249
rect 226 199 618 215
rect 660 249 736 265
rect 660 215 676 249
rect 710 215 736 249
rect 660 199 736 215
rect 778 259 818 282
rect 874 259 914 282
rect 970 259 1010 282
rect 1066 259 1106 282
rect 778 249 1106 259
rect 778 215 802 249
rect 836 215 880 249
rect 914 215 958 249
rect 992 215 1036 249
rect 1070 215 1106 249
rect 226 177 256 199
rect 322 177 352 199
rect 418 177 448 199
rect 514 177 544 199
rect 694 177 724 199
rect 778 198 1106 215
rect 778 177 808 198
rect 880 177 910 198
rect 976 177 1006 198
rect 1076 177 1106 198
rect 1160 265 1200 282
rect 1254 265 1294 282
rect 1348 265 1388 282
rect 1160 249 1418 265
rect 1160 215 1218 249
rect 1252 215 1286 249
rect 1320 215 1364 249
rect 1398 215 1418 249
rect 1160 199 1418 215
rect 1160 177 1190 199
rect 1264 177 1294 199
rect 1360 177 1390 199
rect 120 21 150 47
rect 226 21 256 47
rect 322 21 352 47
rect 418 21 448 47
rect 514 21 544 47
rect 694 21 724 47
rect 778 21 808 47
rect 880 21 910 47
rect 976 21 1006 47
rect 1076 21 1106 47
rect 1160 21 1190 47
rect 1264 21 1294 47
rect 1360 21 1390 47
<< polycont >>
rect 90 215 124 249
rect 292 215 326 249
rect 370 215 404 249
rect 448 215 482 249
rect 676 215 710 249
rect 802 215 836 249
rect 880 215 914 249
rect 958 215 992 249
rect 1036 215 1070 249
rect 1218 215 1252 249
rect 1286 215 1320 249
rect 1364 215 1398 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 19 485 85 493
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 129 485 181 527
rect 129 451 131 485
rect 165 451 181 485
rect 129 435 181 451
rect 236 489 673 493
rect 236 477 437 489
rect 270 455 437 477
rect 471 477 673 489
rect 471 455 635 477
rect 270 443 635 455
rect 669 443 673 477
rect 707 489 783 527
rect 707 455 733 489
rect 767 455 783 489
rect 899 489 975 527
rect 899 455 925 489
rect 959 455 975 489
rect 1019 477 1057 493
rect 19 383 35 417
rect 69 401 85 417
rect 236 409 285 443
rect 411 441 673 443
rect 69 383 202 401
rect 19 357 202 383
rect 270 375 285 409
rect 633 421 673 441
rect 1019 443 1021 477
rect 1055 443 1057 477
rect 1091 489 1167 527
rect 1091 455 1116 489
rect 1150 455 1167 489
rect 1210 477 1247 493
rect 1019 421 1057 443
rect 1244 443 1247 477
rect 1283 489 1359 527
rect 1283 455 1304 489
rect 1338 455 1359 489
rect 1398 477 1448 493
rect 1210 421 1247 443
rect 1432 443 1448 477
rect 1398 421 1448 443
rect 633 415 1448 421
rect 236 359 285 375
rect 336 395 589 407
rect 336 387 533 395
rect 23 249 134 323
rect 23 215 90 249
rect 124 215 134 249
rect 90 199 134 215
rect 168 269 202 357
rect 336 353 341 387
rect 375 361 533 387
rect 567 361 589 395
rect 633 381 829 415
rect 863 409 1448 415
rect 863 381 1021 409
rect 633 375 1021 381
rect 1055 375 1398 409
rect 1432 375 1448 409
rect 375 353 589 361
rect 336 341 589 353
rect 336 317 626 341
rect 168 249 524 269
rect 168 215 292 249
rect 326 215 370 249
rect 404 215 448 249
rect 482 215 524 249
rect 168 207 524 215
rect 168 159 231 207
rect 564 179 626 317
rect 660 296 1424 341
rect 660 249 739 296
rect 660 215 676 249
rect 710 215 739 249
rect 660 213 739 215
rect 773 249 1088 262
rect 773 215 802 249
rect 836 215 880 249
rect 914 215 958 249
rect 992 215 1036 249
rect 1070 215 1088 249
rect 1145 249 1424 296
rect 1145 215 1218 249
rect 1252 215 1286 249
rect 1320 215 1364 249
rect 1398 215 1424 249
rect 773 213 1088 215
rect 564 173 1077 179
rect 18 157 231 159
rect 18 123 39 157
rect 73 123 231 157
rect 275 169 1077 173
rect 275 135 469 169
rect 503 139 835 169
rect 503 135 505 139
rect 711 135 835 139
rect 869 135 1027 169
rect 1061 135 1077 169
rect 1121 164 1365 181
rect 1121 147 1315 164
rect 275 124 505 135
rect 18 89 89 123
rect 275 90 277 124
rect 311 123 505 124
rect 311 90 313 123
rect 18 55 39 89
rect 73 55 89 89
rect 18 51 89 55
rect 154 55 173 89
rect 207 55 231 89
rect 275 74 313 90
rect 467 101 505 123
rect 154 17 231 55
rect 357 55 373 89
rect 407 55 433 89
rect 357 17 433 55
rect 467 67 469 101
rect 503 67 505 101
rect 467 51 505 67
rect 549 89 677 105
rect 1121 101 1173 147
rect 1289 130 1315 147
rect 1349 130 1365 164
rect 549 55 565 89
rect 599 55 643 89
rect 549 17 677 55
rect 713 67 734 101
rect 768 67 931 101
rect 965 89 1173 101
rect 965 67 1116 89
rect 713 55 1116 67
rect 1150 55 1173 89
rect 713 51 1173 55
rect 1217 97 1255 113
rect 1217 63 1219 97
rect 1253 63 1255 97
rect 1217 17 1255 63
rect 1289 96 1365 130
rect 1289 62 1315 96
rect 1349 62 1365 96
rect 1289 51 1365 62
rect 1400 161 1448 177
rect 1434 127 1448 161
rect 1400 93 1448 127
rect 1434 59 1448 93
rect 1400 17 1448 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel locali s 484 357 518 391 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 942 221 976 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 35 289 69 323 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 1145 215 1424 296 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel locali s 660 296 1424 341 1 A2
port 2 nsew signal input
rlabel locali s 660 213 739 296 1 A2
port 2 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_END 189670
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 179800
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
