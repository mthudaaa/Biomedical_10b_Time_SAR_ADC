magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 453 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 267 47 297 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
<< ndiff >>
rect 27 127 89 177
rect 27 93 35 127
rect 69 93 89 127
rect 27 47 89 93
rect 119 95 183 177
rect 119 61 129 95
rect 163 61 183 95
rect 119 47 183 61
rect 213 127 267 177
rect 213 93 223 127
rect 257 93 267 127
rect 213 47 267 93
rect 297 95 427 177
rect 297 61 317 95
rect 351 61 385 95
rect 419 61 427 95
rect 297 47 427 61
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 297 175 497
rect 211 297 269 497
rect 305 485 427 497
rect 305 383 317 485
rect 419 383 427 485
rect 305 297 427 383
<< ndiffc >>
rect 35 93 69 127
rect 129 61 163 95
rect 223 93 257 127
rect 317 61 351 95
rect 385 61 419 95
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 317 383 419 485
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 25 249 119 265
rect 25 215 35 249
rect 69 215 119 249
rect 25 199 119 215
rect 161 249 225 265
rect 161 215 171 249
rect 205 215 225 249
rect 161 199 225 215
rect 267 249 393 265
rect 267 215 349 249
rect 383 215 393 249
rect 267 199 393 215
rect 89 177 119 199
rect 183 177 213 199
rect 267 177 297 199
rect 89 21 119 47
rect 183 21 213 47
rect 267 21 297 47
<< polycont >>
rect 35 215 69 249
rect 171 215 205 249
rect 349 215 383 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 18 485 283 490
rect 18 451 35 485
rect 69 456 283 485
rect 69 451 85 456
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 18 349 85 383
rect 18 315 35 349
rect 69 315 85 349
rect 18 299 85 315
rect 119 265 176 401
rect 18 249 85 265
rect 18 215 35 249
rect 69 215 85 249
rect 18 199 85 215
rect 119 249 215 265
rect 119 215 171 249
rect 205 215 215 249
rect 119 199 215 215
rect 249 165 283 456
rect 317 485 435 527
rect 419 383 435 485
rect 317 367 435 383
rect 18 131 283 165
rect 348 249 441 333
rect 348 215 349 249
rect 383 215 441 249
rect 348 131 441 215
rect 18 127 69 131
rect 18 93 35 127
rect 223 127 257 131
rect 18 77 69 93
rect 103 95 179 97
rect 103 61 129 95
rect 163 61 179 95
rect 223 77 257 93
rect 291 95 435 97
rect 103 17 179 61
rect 291 61 317 95
rect 351 61 385 95
rect 419 61 435 95
rect 291 17 435 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 30 425 64 459 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 392 153 426 187 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 132 289 166 323 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor3_1
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 1722966
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1718370
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
