magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 599 157 795 203
rect 1 21 795 157
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 131
rect 277 47 307 131
rect 349 47 379 131
rect 479 47 509 131
rect 580 47 610 131
rect 687 47 717 177
<< scpmoshvt >>
rect 81 413 117 497
rect 177 413 213 497
rect 299 413 335 497
rect 471 413 507 497
rect 572 413 608 497
rect 679 297 715 497
<< ndiff >>
rect 625 131 687 177
rect 27 101 89 131
rect 27 67 35 101
rect 69 67 89 101
rect 27 47 89 67
rect 119 93 171 131
rect 119 59 129 93
rect 163 59 171 93
rect 119 47 171 59
rect 225 101 277 131
rect 225 67 233 101
rect 267 67 277 101
rect 225 47 277 67
rect 307 47 349 131
rect 379 47 479 131
rect 509 47 580 131
rect 610 93 687 131
rect 610 59 620 93
rect 654 59 687 93
rect 610 47 687 59
rect 717 161 769 177
rect 717 127 727 161
rect 761 127 769 161
rect 717 93 769 127
rect 717 59 727 93
rect 761 59 769 93
rect 717 47 769 59
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 413 81 443
rect 117 485 177 497
rect 117 451 129 485
rect 163 451 177 485
rect 117 413 177 451
rect 213 477 299 497
rect 213 443 240 477
rect 274 443 299 477
rect 213 413 299 443
rect 335 479 471 497
rect 335 445 347 479
rect 381 445 425 479
rect 459 445 471 479
rect 335 413 471 445
rect 507 477 572 497
rect 507 443 526 477
rect 560 443 572 477
rect 507 413 572 443
rect 608 479 679 497
rect 608 445 628 479
rect 662 445 679 479
rect 608 413 679 445
rect 627 297 679 413
rect 715 453 769 497
rect 715 419 727 453
rect 761 419 769 453
rect 715 349 769 419
rect 715 315 727 349
rect 761 315 769 349
rect 715 297 769 315
<< ndiffc >>
rect 35 67 69 101
rect 129 59 163 93
rect 233 67 267 101
rect 620 59 654 93
rect 727 127 761 161
rect 727 59 761 93
<< pdiffc >>
rect 35 443 69 477
rect 129 451 163 485
rect 240 443 274 477
rect 347 445 381 479
rect 425 445 459 479
rect 526 443 560 477
rect 628 445 662 479
rect 727 419 761 453
rect 727 315 761 349
<< poly >>
rect 81 497 117 523
rect 177 497 213 523
rect 299 497 335 523
rect 471 497 507 523
rect 572 497 608 523
rect 679 497 715 523
rect 81 398 117 413
rect 177 398 213 413
rect 299 398 335 413
rect 471 398 507 413
rect 572 398 608 413
rect 79 265 119 398
rect 175 265 215 398
rect 21 249 119 265
rect 21 215 31 249
rect 65 215 119 249
rect 21 199 119 215
rect 161 249 215 265
rect 161 215 171 249
rect 205 215 215 249
rect 297 293 337 398
rect 297 277 379 293
rect 297 243 335 277
rect 369 243 379 277
rect 469 265 509 398
rect 570 265 610 398
rect 679 282 715 297
rect 677 265 717 282
rect 297 227 379 243
rect 161 199 215 215
rect 89 131 119 199
rect 183 176 215 199
rect 183 146 307 176
rect 277 131 307 146
rect 349 131 379 227
rect 455 249 509 265
rect 455 215 465 249
rect 499 215 509 249
rect 455 199 509 215
rect 556 249 610 265
rect 556 215 566 249
rect 600 215 610 249
rect 556 199 610 215
rect 663 249 717 265
rect 663 215 673 249
rect 707 215 717 249
rect 663 199 717 215
rect 479 131 509 199
rect 580 131 610 199
rect 687 177 717 199
rect 89 21 119 47
rect 277 21 307 47
rect 349 21 379 47
rect 479 21 509 47
rect 580 21 610 47
rect 687 21 717 47
<< polycont >>
rect 31 215 65 249
rect 171 215 205 249
rect 335 243 369 277
rect 465 215 499 249
rect 566 215 600 249
rect 673 215 707 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 34 477 69 493
rect 34 443 35 477
rect 34 403 69 443
rect 103 485 179 527
rect 103 451 129 485
rect 163 451 179 485
rect 103 439 179 451
rect 240 477 274 493
rect 331 479 475 527
rect 331 445 347 479
rect 381 445 425 479
rect 459 445 475 479
rect 526 477 560 493
rect 240 409 274 443
rect 612 479 678 527
rect 612 445 628 479
rect 662 445 678 479
rect 727 453 799 493
rect 526 409 560 443
rect 761 419 799 453
rect 34 369 170 403
rect 17 249 90 335
rect 17 215 31 249
rect 65 215 90 249
rect 17 199 90 215
rect 136 265 170 369
rect 240 375 683 409
rect 136 249 205 265
rect 136 215 171 249
rect 136 199 205 215
rect 136 165 170 199
rect 34 131 170 165
rect 34 101 69 131
rect 240 117 274 375
rect 34 67 35 101
rect 228 101 274 117
rect 34 51 69 67
rect 103 59 129 93
rect 163 59 179 93
rect 103 17 179 59
rect 228 67 233 101
rect 267 67 274 101
rect 335 277 431 339
rect 369 243 431 277
rect 335 84 431 243
rect 465 249 523 339
rect 499 215 523 249
rect 465 84 523 215
rect 557 249 615 339
rect 557 215 566 249
rect 600 215 615 249
rect 557 133 615 215
rect 649 265 683 375
rect 727 349 799 419
rect 761 315 799 349
rect 727 299 799 315
rect 649 249 707 265
rect 649 215 673 249
rect 649 199 707 215
rect 745 161 799 299
rect 704 127 727 161
rect 761 127 799 161
rect 704 93 799 127
rect 228 51 274 67
rect 591 59 620 93
rect 654 59 670 93
rect 704 59 727 93
rect 761 59 799 93
rect 591 17 670 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
flabel locali s 470 289 504 323 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 733 85 767 119 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 733 357 767 391 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 733 425 767 459 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 568 221 602 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 568 289 602 323 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 470 85 504 119 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 470 153 504 187 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 376 85 410 119 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 376 153 410 187 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 376 221 410 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 376 289 410 323 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 568 153 602 187 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 470 221 504 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 and4b_1
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 857726
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 849980
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
