
* PEX produced on Sab 26 Okt 2024 02:06:26  CST using ./iic-pex.sh with m=2 and s=1
* NGSPICE file created from delay_element.ext - technology: sky130A
.subckt delay_element_post vdd vip in vin out vss
X0 out a_31_n1616# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=15
X1 a_6375_n1616# vin vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=15
X2 out a_31_n1616# a_6375_n1616# vss sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=15
X3 vss in a_31_n1616# vss sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=15
X4 a_3090_n244# in a_31_n1616# vdd sky130_fd_pr__pfet_01v8_lvt ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=15
X5 vdd vip a_3090_n244# vdd sky130_fd_pr__pfet_01v8_lvt ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=15
C0 a_31_n1616# vin 0.963147f
C1 in vin 1.12606f
C2 a_31_n1616# a_6375_n1616# 0.169373f
C3 vdd vip 7.433569f
C4 vdd a_31_n1616# 6.8485f
C5 vdd in 5.96514f
C6 a_6375_n1616# vin 0.117979f
C7 a_3090_n244# vip 0.41814f
C8 vdd out 0.585541f
C9 vdd vin 0.035251f
C10 a_31_n1616# a_3090_n244# 0.020764f
C11 in a_3090_n244# 0.289501f
C12 a_31_n1616# vip 0.202383f
C13 in vip 1.35686f
C14 in a_31_n1616# 3.37637f
C15 vdd a_3090_n244# 0.977304f
C16 vip vin 0.217406f
C17 a_31_n1616# out 0.479286f
C18 vin vss 11.7144f
C19 out vss 1.23774f
C20 vip vss 4.93206f
C21 in vss 13.5862f
C22 vdd vss 57.480606f
C23 a_6375_n1616# vss 0.825713f $ **FLOATING
C24 a_3090_n244# vss 1.12016f $ **FLOATING
C25 a_31_n1616# vss 15.8812f $ **FLOATING
.ends