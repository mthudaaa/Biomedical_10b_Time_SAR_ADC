magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 1 21 491 203
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 279 47 309 177
rect 377 47 407 177
<< scpmoshvt >>
rect 81 297 117 497
rect 185 297 221 497
rect 281 297 317 497
rect 379 297 415 497
<< ndiff >>
rect 27 95 89 177
rect 27 61 35 95
rect 69 61 89 95
rect 27 47 89 61
rect 119 127 183 177
rect 119 93 129 127
rect 163 93 183 127
rect 119 47 183 93
rect 213 95 279 177
rect 213 61 223 95
rect 257 61 279 95
rect 213 47 279 61
rect 309 127 377 177
rect 309 93 319 127
rect 353 93 377 127
rect 309 47 377 93
rect 407 95 465 177
rect 407 61 417 95
rect 451 61 465 95
rect 407 47 465 61
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 297 185 497
rect 221 297 281 497
rect 317 297 379 497
rect 415 485 469 497
rect 415 451 427 485
rect 461 451 469 485
rect 415 417 469 451
rect 415 383 427 417
rect 461 383 469 417
rect 415 297 469 383
<< ndiffc >>
rect 35 61 69 95
rect 129 93 163 127
rect 223 61 257 95
rect 319 93 353 127
rect 417 61 451 95
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 427 451 461 485
rect 427 383 461 417
<< poly >>
rect 81 497 117 523
rect 185 497 221 523
rect 281 497 317 523
rect 379 497 415 523
rect 81 282 117 297
rect 185 282 221 297
rect 281 282 317 297
rect 379 282 415 297
rect 79 265 119 282
rect 21 249 119 265
rect 21 215 33 249
rect 67 215 119 249
rect 21 199 119 215
rect 89 177 119 199
rect 183 265 223 282
rect 279 265 319 282
rect 377 265 417 282
rect 183 249 237 265
rect 183 215 193 249
rect 227 215 237 249
rect 183 199 237 215
rect 279 249 335 265
rect 279 215 291 249
rect 325 215 335 249
rect 279 199 335 215
rect 377 249 431 265
rect 377 215 387 249
rect 421 215 431 249
rect 377 199 431 215
rect 183 177 213 199
rect 279 177 309 199
rect 377 177 407 199
rect 89 21 119 47
rect 183 21 213 47
rect 279 21 309 47
rect 377 21 407 47
<< polycont >>
rect 33 215 67 249
rect 193 215 227 249
rect 291 215 325 249
rect 387 215 421 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 18 485 85 490
rect 18 451 35 485
rect 69 451 85 485
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 18 349 85 383
rect 18 315 35 349
rect 69 333 85 349
rect 69 315 155 333
rect 18 299 155 315
rect 17 249 67 265
rect 17 215 33 249
rect 17 149 67 215
rect 103 165 155 299
rect 193 249 257 490
rect 227 215 257 249
rect 193 199 257 215
rect 291 249 349 490
rect 427 485 507 527
rect 461 451 507 485
rect 427 417 507 451
rect 461 383 507 417
rect 427 367 507 383
rect 325 215 349 249
rect 291 199 349 215
rect 387 249 441 333
rect 421 215 441 249
rect 103 131 353 165
rect 387 131 441 215
rect 103 127 163 131
rect 17 95 69 115
rect 17 61 35 95
rect 103 93 129 127
rect 319 127 353 131
rect 103 77 163 93
rect 207 95 273 97
rect 17 17 69 61
rect 207 61 223 95
rect 257 61 273 95
rect 319 77 353 93
rect 401 95 504 97
rect 207 17 273 61
rect 401 61 417 95
rect 451 61 504 95
rect 401 17 504 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel locali s 29 153 63 187 0 FreeSans 400 0 0 0 D
port 4 nsew signal input
flabel locali s 207 289 241 323 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 28 221 62 255 0 FreeSans 400 0 0 0 D
port 4 nsew signal input
flabel locali s 30 425 64 459 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 394 153 428 187 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 301 357 335 391 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4_1
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 1768334
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1763454
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
