magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 163 197 203
rect 523 163 725 203
rect 1 67 725 163
rect 30 27 725 67
rect 30 -17 64 27
rect 526 21 725 27
<< scnmos >>
rect 89 93 119 177
rect 287 53 317 137
rect 381 53 411 137
rect 462 53 492 137
rect 617 47 647 177
<< scpmoshvt >>
rect 81 413 117 497
rect 279 311 315 395
rect 373 311 409 395
rect 478 297 514 381
rect 609 297 645 497
<< ndiff >>
rect 27 163 89 177
rect 27 129 35 163
rect 69 129 89 163
rect 27 93 89 129
rect 119 165 171 177
rect 119 131 129 165
rect 163 131 171 165
rect 549 137 617 177
rect 119 93 171 131
rect 230 99 287 137
rect 230 65 238 99
rect 272 65 287 99
rect 230 53 287 65
rect 317 53 381 137
rect 411 53 462 137
rect 492 109 617 137
rect 492 75 571 109
rect 605 75 617 109
rect 492 53 617 75
rect 552 47 617 53
rect 647 119 699 177
rect 647 85 657 119
rect 691 85 699 119
rect 647 47 699 85
<< pdiff >>
rect 27 475 81 497
rect 27 441 35 475
rect 69 441 81 475
rect 27 413 81 441
rect 117 469 171 497
rect 117 435 129 469
rect 163 435 171 469
rect 117 413 171 435
rect 555 485 609 497
rect 555 451 563 485
rect 597 451 609 485
rect 225 369 279 395
rect 225 335 233 369
rect 267 335 279 369
rect 225 311 279 335
rect 315 387 373 395
rect 315 353 327 387
rect 361 353 373 387
rect 315 311 373 353
rect 409 381 461 395
rect 555 381 609 451
rect 409 362 478 381
rect 409 328 431 362
rect 465 328 478 362
rect 409 311 478 328
rect 426 297 478 311
rect 514 297 609 381
rect 645 471 699 497
rect 645 437 657 471
rect 691 437 699 471
rect 645 403 699 437
rect 645 369 657 403
rect 691 369 699 403
rect 645 297 699 369
<< ndiffc >>
rect 35 129 69 163
rect 129 131 163 165
rect 238 65 272 99
rect 571 75 605 109
rect 657 85 691 119
<< pdiffc >>
rect 35 441 69 475
rect 129 435 163 469
rect 563 451 597 485
rect 233 335 267 369
rect 327 353 361 387
rect 431 328 465 362
rect 657 437 691 471
rect 657 369 691 403
<< poly >>
rect 81 497 117 523
rect 371 477 438 500
rect 609 497 645 523
rect 371 443 384 477
rect 418 443 438 477
rect 371 427 438 443
rect 81 398 117 413
rect 79 339 119 398
rect 279 395 315 425
rect 371 421 411 427
rect 373 395 409 421
rect 22 323 119 339
rect 22 289 35 323
rect 69 289 119 323
rect 478 381 514 407
rect 279 296 315 311
rect 373 296 409 311
rect 22 249 119 289
rect 277 265 317 296
rect 22 215 35 249
rect 69 215 119 249
rect 22 199 119 215
rect 243 249 317 265
rect 243 215 253 249
rect 287 215 317 249
rect 371 240 411 296
rect 478 282 514 297
rect 609 282 645 297
rect 476 265 516 282
rect 607 265 647 282
rect 243 199 317 215
rect 89 177 119 199
rect 287 137 317 199
rect 381 137 411 240
rect 462 249 516 265
rect 462 215 472 249
rect 506 215 516 249
rect 462 199 516 215
rect 593 249 647 265
rect 593 215 603 249
rect 637 215 647 249
rect 593 199 647 215
rect 462 137 492 199
rect 617 177 647 199
rect 89 67 119 93
rect 287 27 317 53
rect 381 27 411 53
rect 462 27 492 53
rect 617 21 647 47
<< polycont >>
rect 384 443 418 477
rect 35 289 69 323
rect 35 215 69 249
rect 253 215 287 249
rect 472 215 506 249
rect 603 215 637 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 475 69 527
rect 17 441 35 475
rect 17 425 69 441
rect 129 469 163 493
rect 17 323 85 391
rect 17 289 35 323
rect 69 289 85 323
rect 17 249 85 289
rect 17 215 35 249
rect 69 215 85 249
rect 129 249 163 435
rect 217 426 350 527
rect 301 391 350 426
rect 384 477 499 493
rect 418 443 499 477
rect 384 425 499 443
rect 559 485 602 527
rect 559 451 563 485
rect 597 451 602 485
rect 559 418 602 451
rect 654 471 707 493
rect 654 437 657 471
rect 691 437 707 471
rect 654 403 707 437
rect 217 369 267 388
rect 217 335 233 369
rect 301 387 377 391
rect 301 353 327 387
rect 361 353 377 387
rect 431 362 610 378
rect 217 319 267 335
rect 465 328 610 362
rect 654 369 657 403
rect 691 369 707 403
rect 654 353 707 369
rect 431 319 610 328
rect 217 315 610 319
rect 217 285 637 315
rect 129 215 253 249
rect 287 215 304 249
rect 129 199 304 215
rect 129 181 179 199
rect 17 163 69 181
rect 17 129 35 163
rect 17 17 69 129
rect 103 165 179 181
rect 103 131 129 165
rect 163 131 179 165
rect 103 97 179 131
rect 338 110 389 285
rect 221 99 389 110
rect 221 65 238 99
rect 272 65 389 99
rect 221 57 389 65
rect 456 249 529 251
rect 456 215 472 249
rect 506 215 529 249
rect 456 61 529 215
rect 593 249 637 285
rect 593 215 603 249
rect 593 195 637 215
rect 673 147 707 353
rect 563 109 621 125
rect 563 75 571 109
rect 605 75 621 109
rect 563 17 621 75
rect 655 119 707 147
rect 655 85 657 119
rect 691 85 707 119
rect 655 51 707 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 30 289 64 323 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel locali s 384 425 499 493 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 663 425 697 459 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 473 153 507 187 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel locali s 660 85 694 119 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 30 357 64 391 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 and3b_1
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 814124
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 807718
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
