magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 23 201 1737 203
rect 23 23 2078 201
rect 23 21 513 23
rect 1001 21 1213 23
rect 1652 21 2078 23
rect 29 -17 63 21
<< scnmos >>
rect 101 47 131 177
rect 195 47 225 177
rect 291 47 321 177
rect 385 47 415 177
rect 502 93 532 177
rect 745 49 775 177
rect 851 49 881 177
rect 1095 47 1125 177
rect 1301 49 1331 177
rect 1462 49 1492 133
rect 1621 49 1651 177
rect 1761 47 1791 167
rect 1871 47 1901 175
rect 1965 47 1995 175
<< scpmoshvt >>
rect 103 297 139 497
rect 197 297 233 497
rect 297 297 333 497
rect 391 297 427 497
rect 504 297 540 425
rect 724 325 760 493
rect 831 297 867 465
rect 1053 297 1089 497
rect 1293 297 1329 465
rect 1454 297 1490 425
rect 1639 329 1675 457
rect 1752 329 1788 497
rect 1863 297 1899 497
rect 1957 297 1993 497
<< ndiff >>
rect 49 129 101 177
rect 49 95 57 129
rect 91 95 101 129
rect 49 47 101 95
rect 131 129 195 177
rect 131 95 151 129
rect 185 95 195 129
rect 131 47 195 95
rect 225 129 291 177
rect 225 95 245 129
rect 279 95 291 129
rect 225 47 291 95
rect 321 129 385 177
rect 321 95 341 129
rect 375 95 385 129
rect 321 47 385 95
rect 415 93 502 177
rect 532 169 627 177
rect 532 135 581 169
rect 615 135 627 169
rect 532 93 627 135
rect 681 165 745 177
rect 681 131 691 165
rect 725 131 745 165
rect 415 89 487 93
rect 415 55 435 89
rect 469 55 487 89
rect 415 47 487 55
rect 681 49 745 131
rect 775 91 851 177
rect 775 57 787 91
rect 821 57 851 91
rect 775 49 851 57
rect 881 91 943 177
rect 881 57 897 91
rect 931 57 943 91
rect 881 49 943 57
rect 1027 157 1095 177
rect 1027 123 1041 157
rect 1075 123 1095 157
rect 1027 89 1095 123
rect 1027 55 1041 89
rect 1075 55 1095 89
rect 1027 47 1095 55
rect 1125 165 1187 177
rect 1125 131 1145 165
rect 1179 131 1187 165
rect 1125 47 1187 131
rect 1241 97 1301 177
rect 1241 63 1254 97
rect 1288 63 1301 97
rect 1241 49 1301 63
rect 1331 133 1431 177
rect 1517 169 1621 177
rect 1517 135 1563 169
rect 1597 135 1621 169
rect 1517 133 1621 135
rect 1331 126 1462 133
rect 1331 92 1341 126
rect 1375 92 1462 126
rect 1331 49 1462 92
rect 1492 49 1621 133
rect 1651 167 1711 177
rect 1811 167 1871 175
rect 1651 93 1761 167
rect 1651 59 1673 93
rect 1707 59 1761 93
rect 1651 49 1761 59
rect 1678 47 1761 49
rect 1791 142 1871 167
rect 1791 108 1817 142
rect 1851 108 1871 142
rect 1791 47 1871 108
rect 1901 97 1965 175
rect 1901 63 1911 97
rect 1945 63 1965 97
rect 1901 47 1965 63
rect 1995 101 2052 175
rect 1995 67 2005 101
rect 2039 67 2052 101
rect 1995 47 2052 67
<< pdiff >>
rect 49 485 103 497
rect 49 451 57 485
rect 91 451 103 485
rect 49 417 103 451
rect 49 383 57 417
rect 91 383 103 417
rect 49 349 103 383
rect 49 315 57 349
rect 91 315 103 349
rect 49 297 103 315
rect 139 485 197 497
rect 139 451 151 485
rect 185 451 197 485
rect 139 417 197 451
rect 139 383 151 417
rect 185 383 197 417
rect 139 349 197 383
rect 139 315 151 349
rect 185 315 197 349
rect 139 297 197 315
rect 233 485 297 497
rect 233 451 245 485
rect 279 451 297 485
rect 233 417 297 451
rect 233 383 245 417
rect 279 383 297 417
rect 233 349 297 383
rect 233 315 245 349
rect 279 315 297 349
rect 233 297 297 315
rect 333 477 391 497
rect 333 443 345 477
rect 379 443 391 477
rect 333 409 391 443
rect 333 375 345 409
rect 379 375 391 409
rect 333 341 391 375
rect 333 307 345 341
rect 379 307 391 341
rect 333 297 391 307
rect 427 477 487 497
rect 427 443 440 477
rect 474 443 487 477
rect 427 425 487 443
rect 427 297 504 425
rect 540 341 598 425
rect 540 307 552 341
rect 586 307 598 341
rect 657 413 724 493
rect 657 379 678 413
rect 712 379 724 413
rect 657 325 724 379
rect 760 481 814 493
rect 760 447 772 481
rect 806 465 814 481
rect 999 481 1053 497
rect 806 447 831 465
rect 760 325 831 447
rect 540 297 598 307
rect 779 297 831 325
rect 867 423 945 465
rect 999 447 1007 481
rect 1041 447 1053 481
rect 999 435 1053 447
rect 867 339 946 423
rect 867 305 900 339
rect 934 305 946 339
rect 867 297 946 305
rect 1000 297 1053 435
rect 1089 343 1153 497
rect 1692 489 1752 497
rect 1089 309 1101 343
rect 1135 309 1153 343
rect 1089 297 1153 309
rect 1207 405 1293 465
rect 1207 371 1215 405
rect 1249 371 1293 405
rect 1207 297 1293 371
rect 1329 425 1430 465
rect 1692 457 1704 489
rect 1552 425 1639 457
rect 1329 409 1454 425
rect 1329 375 1381 409
rect 1415 375 1454 409
rect 1329 341 1454 375
rect 1329 307 1381 341
rect 1415 307 1454 341
rect 1329 297 1454 307
rect 1490 421 1639 425
rect 1490 387 1593 421
rect 1627 387 1639 421
rect 1490 329 1639 387
rect 1675 455 1704 457
rect 1738 455 1752 489
rect 1675 329 1752 455
rect 1788 341 1863 497
rect 1788 329 1817 341
rect 1490 297 1587 329
rect 1805 307 1817 329
rect 1851 307 1863 341
rect 1805 297 1863 307
rect 1899 489 1957 497
rect 1899 455 1911 489
rect 1945 455 1957 489
rect 1899 297 1957 455
rect 1993 477 2052 497
rect 1993 443 2006 477
rect 2040 443 2052 477
rect 1993 409 2052 443
rect 1993 375 2006 409
rect 2040 375 2052 409
rect 1993 297 2052 375
<< ndiffc >>
rect 57 95 91 129
rect 151 95 185 129
rect 245 95 279 129
rect 341 95 375 129
rect 581 135 615 169
rect 691 131 725 165
rect 435 55 469 89
rect 787 57 821 91
rect 897 57 931 91
rect 1041 123 1075 157
rect 1041 55 1075 89
rect 1145 131 1179 165
rect 1254 63 1288 97
rect 1563 135 1597 169
rect 1341 92 1375 126
rect 1673 59 1707 93
rect 1817 108 1851 142
rect 1911 63 1945 97
rect 2005 67 2039 101
<< pdiffc >>
rect 57 451 91 485
rect 57 383 91 417
rect 57 315 91 349
rect 151 451 185 485
rect 151 383 185 417
rect 151 315 185 349
rect 245 451 279 485
rect 245 383 279 417
rect 245 315 279 349
rect 345 443 379 477
rect 345 375 379 409
rect 345 307 379 341
rect 440 443 474 477
rect 552 307 586 341
rect 678 379 712 413
rect 772 447 806 481
rect 1007 447 1041 481
rect 900 305 934 339
rect 1101 309 1135 343
rect 1215 371 1249 405
rect 1381 375 1415 409
rect 1381 307 1415 341
rect 1593 387 1627 421
rect 1704 455 1738 489
rect 1817 307 1851 341
rect 1911 455 1945 489
rect 2006 443 2040 477
rect 2006 375 2040 409
<< poly >>
rect 103 497 139 523
rect 197 497 233 523
rect 297 497 333 523
rect 391 497 427 523
rect 724 493 760 519
rect 502 451 542 483
rect 504 425 540 451
rect 831 465 867 504
rect 1053 497 1089 523
rect 724 310 760 325
rect 103 282 139 297
rect 197 282 233 297
rect 297 282 333 297
rect 391 282 427 297
rect 504 282 540 297
rect 101 265 141 282
rect 195 265 235 282
rect 295 265 335 282
rect 389 265 429 282
rect 502 265 542 282
rect 722 271 762 310
rect 1291 493 1677 523
rect 1752 497 1788 523
rect 1863 497 1899 523
rect 1957 497 1993 523
rect 1291 491 1331 493
rect 1293 465 1329 491
rect 1637 483 1677 493
rect 1639 457 1675 483
rect 1454 425 1490 451
rect 1639 314 1675 329
rect 1752 314 1788 329
rect 831 282 867 297
rect 1053 282 1089 297
rect 1293 282 1329 297
rect 1454 282 1490 297
rect 722 265 775 271
rect 829 265 869 282
rect 101 249 460 265
rect 101 215 406 249
rect 440 215 460 249
rect 101 199 460 215
rect 502 249 775 265
rect 502 215 692 249
rect 726 215 775 249
rect 502 199 775 215
rect 817 249 881 265
rect 817 215 827 249
rect 861 215 881 249
rect 1051 247 1091 282
rect 1291 247 1331 282
rect 1452 265 1492 282
rect 1637 265 1677 314
rect 1051 217 1331 247
rect 817 199 881 215
rect 101 177 131 199
rect 195 177 225 199
rect 291 177 321 199
rect 385 177 415 199
rect 502 177 532 199
rect 745 177 775 199
rect 851 177 881 199
rect 1095 177 1125 217
rect 1301 177 1331 217
rect 1373 249 1492 265
rect 1373 215 1383 249
rect 1417 215 1492 249
rect 1373 199 1492 215
rect 502 67 532 93
rect 101 21 131 47
rect 195 21 225 47
rect 291 21 321 47
rect 385 21 415 47
rect 745 21 775 49
rect 851 21 881 49
rect 1462 133 1492 199
rect 1621 249 1685 265
rect 1750 256 1790 314
rect 1863 282 1899 297
rect 1957 282 1993 297
rect 1861 265 1901 282
rect 1955 265 1995 282
rect 1750 255 1791 256
rect 1621 215 1631 249
rect 1665 215 1685 249
rect 1621 199 1685 215
rect 1727 239 1791 255
rect 1727 205 1737 239
rect 1771 205 1791 239
rect 1621 177 1651 199
rect 1727 189 1791 205
rect 1833 249 1901 265
rect 1833 215 1843 249
rect 1877 215 1901 249
rect 1833 199 1901 215
rect 1943 249 2007 265
rect 1943 215 1953 249
rect 1987 215 2007 249
rect 1943 199 2007 215
rect 1761 167 1791 189
rect 1871 175 1901 199
rect 1965 175 1995 199
rect 1095 21 1125 47
rect 1301 21 1331 49
rect 1462 23 1492 49
rect 1621 21 1651 49
rect 1761 21 1791 47
rect 1871 21 1901 47
rect 1965 21 1995 47
<< polycont >>
rect 406 215 440 249
rect 692 215 726 249
rect 827 215 861 249
rect 1383 215 1417 249
rect 1631 215 1665 249
rect 1737 205 1771 239
rect 1843 215 1877 249
rect 1953 215 1987 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 57 485 91 527
rect 245 485 279 527
rect 57 417 91 451
rect 57 349 91 383
rect 57 298 91 315
rect 125 451 151 485
rect 185 451 201 485
rect 125 417 201 451
rect 125 383 151 417
rect 185 383 201 417
rect 125 349 201 383
rect 125 315 151 349
rect 185 315 201 349
rect 125 265 201 315
rect 245 417 279 451
rect 245 349 279 383
rect 245 299 279 315
rect 313 477 379 493
rect 313 443 345 477
rect 413 477 490 527
rect 991 481 1057 527
rect 1885 489 1962 527
rect 413 443 440 477
rect 474 443 490 477
rect 526 447 772 481
rect 806 447 840 481
rect 991 447 1007 481
rect 1041 447 1057 481
rect 1144 455 1704 489
rect 1738 455 1803 489
rect 1885 455 1911 489
rect 1945 455 1962 489
rect 2006 477 2065 493
rect 313 409 379 443
rect 526 409 570 447
rect 1144 413 1178 455
rect 313 375 345 409
rect 313 341 379 375
rect 313 307 345 341
rect 313 288 379 307
rect 413 375 570 409
rect 638 379 678 413
rect 712 379 1178 413
rect 1215 405 1249 421
rect 313 265 372 288
rect 413 265 457 375
rect 503 307 552 341
rect 586 307 840 341
rect 125 199 372 265
rect 406 249 457 265
rect 440 215 457 249
rect 406 199 457 215
rect 57 129 91 147
rect 57 17 91 95
rect 125 129 185 199
rect 313 185 372 199
rect 125 95 151 129
rect 125 75 185 95
rect 245 129 279 147
rect 245 17 279 95
rect 313 129 375 185
rect 412 173 457 199
rect 412 139 547 173
rect 313 95 341 129
rect 313 70 375 95
rect 409 89 469 105
rect 409 55 435 89
rect 409 17 469 55
rect 503 85 547 139
rect 581 169 615 307
rect 806 265 840 307
rect 884 305 900 339
rect 934 323 961 339
rect 905 289 927 305
rect 905 275 961 289
rect 649 249 772 265
rect 649 215 692 249
rect 726 215 772 249
rect 806 249 871 265
rect 806 215 827 249
rect 861 215 871 249
rect 806 199 871 215
rect 581 119 615 135
rect 675 165 751 181
rect 675 131 691 165
rect 725 159 751 165
rect 905 159 939 275
rect 995 241 1029 379
rect 1075 309 1101 343
rect 1135 309 1179 343
rect 1075 289 1179 309
rect 725 131 939 159
rect 675 125 939 131
rect 973 207 1029 241
rect 973 91 1007 207
rect 1121 187 1179 289
rect 740 85 787 91
rect 503 57 787 85
rect 821 57 837 91
rect 881 57 897 91
rect 931 57 1007 91
rect 1041 157 1075 173
rect 1041 89 1075 123
rect 503 51 837 57
rect 1155 165 1179 187
rect 1121 131 1145 153
rect 1121 83 1179 131
rect 1215 119 1249 371
rect 1283 165 1317 455
rect 2040 443 2065 477
rect 2006 421 2065 443
rect 1363 375 1381 409
rect 1415 375 1446 409
rect 1363 341 1446 375
rect 1363 307 1381 341
rect 1415 323 1446 341
rect 1563 387 1593 421
rect 1627 409 2065 421
rect 1627 387 2006 409
rect 1415 307 1417 323
rect 1363 289 1417 307
rect 1451 289 1529 323
rect 1366 249 1451 254
rect 1366 215 1383 249
rect 1417 215 1451 249
rect 1366 199 1451 215
rect 1409 187 1451 199
rect 1283 131 1375 165
rect 1341 126 1375 131
rect 1409 153 1417 187
rect 1409 126 1451 153
rect 1249 85 1254 97
rect 1041 17 1075 55
rect 1215 63 1254 85
rect 1288 63 1304 97
rect 1341 64 1375 92
rect 1495 85 1529 289
rect 1563 169 1597 387
rect 1958 375 2006 387
rect 2040 375 2065 409
rect 1631 289 1757 323
rect 1801 307 1817 341
rect 1851 307 1975 341
rect 1801 299 1975 307
rect 1631 249 1675 289
rect 1941 265 1975 299
rect 1665 215 1675 249
rect 1631 199 1675 215
rect 1709 239 1771 255
rect 1709 205 1737 239
rect 1815 249 1907 265
rect 1815 215 1843 249
rect 1877 215 1907 249
rect 1941 249 1997 265
rect 1941 215 1953 249
rect 1987 215 1997 249
rect 1709 189 1771 205
rect 1941 199 1997 215
rect 1709 187 1750 189
rect 1709 153 1713 187
rect 1747 153 1750 187
rect 1941 181 1975 199
rect 1709 146 1750 153
rect 1817 150 1975 181
rect 1809 147 1975 150
rect 1563 119 1597 135
rect 1809 142 1867 147
rect 1809 119 1817 142
rect 1631 85 1673 93
rect 1215 53 1304 63
rect 1495 59 1673 85
rect 1707 59 1734 93
rect 1809 85 1815 119
rect 1851 108 1867 142
rect 2031 117 2065 375
rect 1849 85 1867 108
rect 1809 59 1867 85
rect 1911 97 1945 113
rect 1495 51 1734 59
rect 1911 17 1945 63
rect 2005 101 2065 117
rect 2039 67 2065 101
rect 2005 51 2065 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 927 305 934 323
rect 934 305 961 323
rect 927 289 961 305
rect 1121 165 1155 187
rect 1121 153 1145 165
rect 1145 153 1155 165
rect 1417 289 1451 323
rect 1215 85 1249 119
rect 1417 153 1451 187
rect 1713 153 1747 187
rect 1815 108 1817 119
rect 1817 108 1849 119
rect 1815 85 1849 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 915 323 973 329
rect 915 289 927 323
rect 961 320 973 323
rect 1405 323 1463 329
rect 1405 320 1417 323
rect 961 292 1417 320
rect 961 289 973 292
rect 915 283 973 289
rect 1405 289 1417 292
rect 1451 289 1463 323
rect 1405 283 1463 289
rect 1109 187 1167 193
rect 1109 153 1121 187
rect 1155 184 1167 187
rect 1405 187 1463 193
rect 1405 184 1417 187
rect 1155 156 1417 184
rect 1155 153 1167 156
rect 1109 147 1167 153
rect 1405 153 1417 156
rect 1451 184 1463 187
rect 1701 187 1759 193
rect 1701 184 1713 187
rect 1451 156 1713 184
rect 1451 153 1463 156
rect 1405 147 1463 153
rect 1701 153 1713 156
rect 1747 153 1759 187
rect 1701 147 1759 153
rect 1203 119 1263 125
rect 1203 85 1215 119
rect 1249 116 1263 119
rect 1803 119 1861 125
rect 1803 116 1815 119
rect 1249 88 1815 116
rect 1249 85 1263 88
rect 1203 79 1263 85
rect 1803 85 1815 88
rect 1849 85 1861 119
rect 1803 79 1861 85
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< labels >>
flabel locali s 319 357 353 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1689 289 1723 323 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1815 215 1907 265 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 hkscl5hdv1_xnor3_1
flabel comment s 0 544 0 544 3 FreeSans 200 0 0 0 HHNEC
<< properties >>
string FIXED_BBOX 0 0 2116 544
string GDS_END 2814750
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 2800828
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
