magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 1 21 2203 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 458 47 488 177
rect 552 47 582 177
rect 646 47 676 177
rect 750 47 780 177
rect 834 47 864 177
rect 928 47 958 177
rect 1022 47 1052 177
rect 1148 47 1178 177
rect 1314 47 1344 177
rect 1408 47 1438 177
rect 1502 47 1532 177
rect 1606 47 1636 177
rect 1794 47 1824 177
rect 1888 47 1918 177
rect 1982 47 2012 177
rect 2085 47 2115 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 460 297 496 497
rect 554 297 590 497
rect 648 297 684 497
rect 742 297 778 497
rect 940 297 976 497
rect 1034 297 1070 497
rect 1128 297 1164 497
rect 1222 297 1258 497
rect 1316 297 1352 497
rect 1410 297 1446 497
rect 1504 297 1540 497
rect 1598 297 1634 497
rect 1796 297 1832 497
rect 1890 297 1926 497
rect 1984 297 2020 497
rect 2087 297 2123 497
<< ndiff >>
rect 27 161 89 177
rect 27 127 35 161
rect 69 127 89 161
rect 27 93 89 127
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 165 183 177
rect 119 131 129 165
rect 163 131 183 165
rect 119 47 183 131
rect 213 93 277 177
rect 213 59 223 93
rect 257 59 277 93
rect 213 47 277 59
rect 307 165 371 177
rect 307 131 317 165
rect 351 131 371 165
rect 307 47 371 131
rect 401 93 458 177
rect 401 59 411 93
rect 445 59 458 93
rect 401 47 458 59
rect 488 165 552 177
rect 488 131 508 165
rect 542 131 552 165
rect 488 47 552 131
rect 582 93 646 177
rect 582 59 602 93
rect 636 59 646 93
rect 582 47 646 59
rect 676 165 750 177
rect 676 131 696 165
rect 730 131 750 165
rect 676 47 750 131
rect 780 165 834 177
rect 780 131 790 165
rect 824 131 834 165
rect 780 93 834 131
rect 780 59 790 93
rect 824 59 834 93
rect 780 47 834 59
rect 864 93 928 177
rect 864 59 884 93
rect 918 59 928 93
rect 864 47 928 59
rect 958 165 1022 177
rect 958 131 978 165
rect 1012 131 1022 165
rect 958 93 1022 131
rect 958 59 978 93
rect 1012 59 1022 93
rect 958 47 1022 59
rect 1052 93 1148 177
rect 1052 59 1088 93
rect 1122 59 1148 93
rect 1052 47 1148 59
rect 1178 165 1314 177
rect 1178 131 1198 165
rect 1232 131 1266 165
rect 1300 131 1314 165
rect 1178 93 1314 131
rect 1178 59 1198 93
rect 1232 59 1266 93
rect 1300 59 1314 93
rect 1178 47 1314 59
rect 1344 93 1408 177
rect 1344 59 1364 93
rect 1398 59 1408 93
rect 1344 47 1408 59
rect 1438 165 1502 177
rect 1438 131 1458 165
rect 1492 131 1502 165
rect 1438 93 1502 131
rect 1438 59 1458 93
rect 1492 59 1502 93
rect 1438 47 1502 59
rect 1532 93 1606 177
rect 1532 59 1552 93
rect 1586 59 1606 93
rect 1532 47 1606 59
rect 1636 165 1794 177
rect 1636 131 1646 165
rect 1680 131 1718 165
rect 1752 131 1794 165
rect 1636 93 1794 131
rect 1636 59 1646 93
rect 1680 59 1718 93
rect 1752 59 1794 93
rect 1636 47 1794 59
rect 1824 93 1888 177
rect 1824 59 1844 93
rect 1878 59 1888 93
rect 1824 47 1888 59
rect 1918 165 1982 177
rect 1918 131 1938 165
rect 1972 131 1982 165
rect 1918 93 1982 131
rect 1918 59 1938 93
rect 1972 59 1982 93
rect 1918 47 1982 59
rect 2012 93 2085 177
rect 2012 59 2041 93
rect 2075 59 2085 93
rect 2012 47 2085 59
rect 2115 165 2177 177
rect 2115 131 2135 165
rect 2169 131 2177 165
rect 2115 93 2177 131
rect 2115 59 2135 93
rect 2169 59 2177 93
rect 2115 47 2177 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 417 175 497
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 417 363 497
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 451 460 497
rect 399 417 414 451
rect 448 417 460 451
rect 399 297 460 417
rect 496 485 554 497
rect 496 451 508 485
rect 542 451 554 485
rect 496 297 554 451
rect 590 469 648 497
rect 590 435 602 469
rect 636 435 648 469
rect 590 401 648 435
rect 590 367 602 401
rect 636 367 648 401
rect 590 297 648 367
rect 684 485 742 497
rect 684 451 696 485
rect 730 451 742 485
rect 684 297 742 451
rect 778 469 832 497
rect 778 435 790 469
rect 824 435 832 469
rect 778 401 832 435
rect 778 367 790 401
rect 824 367 832 401
rect 778 297 832 367
rect 886 485 940 497
rect 886 451 894 485
rect 928 451 940 485
rect 886 417 940 451
rect 886 383 894 417
rect 928 383 940 417
rect 886 297 940 383
rect 976 417 1034 497
rect 976 383 988 417
rect 1022 383 1034 417
rect 976 349 1034 383
rect 976 315 988 349
rect 1022 315 1034 349
rect 976 297 1034 315
rect 1070 485 1128 497
rect 1070 451 1082 485
rect 1116 451 1128 485
rect 1070 417 1128 451
rect 1070 383 1082 417
rect 1116 383 1128 417
rect 1070 297 1128 383
rect 1164 417 1222 497
rect 1164 383 1176 417
rect 1210 383 1222 417
rect 1164 349 1222 383
rect 1164 315 1176 349
rect 1210 315 1222 349
rect 1164 297 1222 315
rect 1258 485 1316 497
rect 1258 451 1270 485
rect 1304 451 1316 485
rect 1258 417 1316 451
rect 1258 383 1270 417
rect 1304 383 1316 417
rect 1258 297 1316 383
rect 1352 417 1410 497
rect 1352 383 1364 417
rect 1398 383 1410 417
rect 1352 349 1410 383
rect 1352 315 1364 349
rect 1398 315 1410 349
rect 1352 297 1410 315
rect 1446 485 1504 497
rect 1446 451 1458 485
rect 1492 451 1504 485
rect 1446 417 1504 451
rect 1446 383 1458 417
rect 1492 383 1504 417
rect 1446 297 1504 383
rect 1540 417 1598 497
rect 1540 383 1552 417
rect 1586 383 1598 417
rect 1540 349 1598 383
rect 1540 315 1552 349
rect 1586 315 1598 349
rect 1540 297 1598 315
rect 1634 485 1688 497
rect 1634 451 1646 485
rect 1680 451 1688 485
rect 1634 417 1688 451
rect 1634 383 1646 417
rect 1680 383 1688 417
rect 1634 297 1688 383
rect 1742 485 1796 497
rect 1742 451 1750 485
rect 1784 451 1796 485
rect 1742 417 1796 451
rect 1742 383 1750 417
rect 1784 383 1796 417
rect 1742 297 1796 383
rect 1832 485 1890 497
rect 1832 451 1844 485
rect 1878 451 1890 485
rect 1832 417 1890 451
rect 1832 383 1844 417
rect 1878 383 1890 417
rect 1832 349 1890 383
rect 1832 315 1844 349
rect 1878 315 1890 349
rect 1832 297 1890 315
rect 1926 485 1984 497
rect 1926 451 1938 485
rect 1972 451 1984 485
rect 1926 417 1984 451
rect 1926 383 1938 417
rect 1972 383 1984 417
rect 1926 297 1984 383
rect 2020 485 2087 497
rect 2020 451 2032 485
rect 2066 451 2087 485
rect 2020 417 2087 451
rect 2020 383 2032 417
rect 2066 383 2087 417
rect 2020 349 2087 383
rect 2020 315 2032 349
rect 2066 315 2087 349
rect 2020 297 2087 315
rect 2123 485 2177 497
rect 2123 451 2135 485
rect 2169 451 2177 485
rect 2123 417 2177 451
rect 2123 383 2135 417
rect 2169 383 2177 417
rect 2123 349 2177 383
rect 2123 315 2135 349
rect 2169 315 2177 349
rect 2123 297 2177 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 131 163 165
rect 223 59 257 93
rect 317 131 351 165
rect 411 59 445 93
rect 508 131 542 165
rect 602 59 636 93
rect 696 131 730 165
rect 790 131 824 165
rect 790 59 824 93
rect 884 59 918 93
rect 978 131 1012 165
rect 978 59 1012 93
rect 1088 59 1122 93
rect 1198 131 1232 165
rect 1266 131 1300 165
rect 1198 59 1232 93
rect 1266 59 1300 93
rect 1364 59 1398 93
rect 1458 131 1492 165
rect 1458 59 1492 93
rect 1552 59 1586 93
rect 1646 131 1680 165
rect 1718 131 1752 165
rect 1646 59 1680 93
rect 1718 59 1752 93
rect 1844 59 1878 93
rect 1938 131 1972 165
rect 1938 59 1972 93
rect 2041 59 2075 93
rect 2135 131 2169 165
rect 2135 59 2169 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 383 351 417
rect 317 315 351 349
rect 414 417 448 451
rect 508 451 542 485
rect 602 435 636 469
rect 602 367 636 401
rect 696 451 730 485
rect 790 435 824 469
rect 790 367 824 401
rect 894 451 928 485
rect 894 383 928 417
rect 988 383 1022 417
rect 988 315 1022 349
rect 1082 451 1116 485
rect 1082 383 1116 417
rect 1176 383 1210 417
rect 1176 315 1210 349
rect 1270 451 1304 485
rect 1270 383 1304 417
rect 1364 383 1398 417
rect 1364 315 1398 349
rect 1458 451 1492 485
rect 1458 383 1492 417
rect 1552 383 1586 417
rect 1552 315 1586 349
rect 1646 451 1680 485
rect 1646 383 1680 417
rect 1750 451 1784 485
rect 1750 383 1784 417
rect 1844 451 1878 485
rect 1844 383 1878 417
rect 1844 315 1878 349
rect 1938 451 1972 485
rect 1938 383 1972 417
rect 2032 451 2066 485
rect 2032 383 2066 417
rect 2032 315 2066 349
rect 2135 451 2169 485
rect 2135 383 2169 417
rect 2135 315 2169 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 460 497 496 523
rect 554 497 590 523
rect 648 497 684 523
rect 742 497 778 523
rect 940 497 976 523
rect 1034 497 1070 523
rect 1128 497 1164 523
rect 1222 497 1258 523
rect 1316 497 1352 523
rect 1410 497 1446 523
rect 1504 497 1540 523
rect 1598 497 1634 523
rect 1796 497 1832 523
rect 1890 497 1926 523
rect 1984 497 2020 523
rect 2087 497 2123 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 460 282 496 297
rect 554 282 590 297
rect 648 282 684 297
rect 742 282 778 297
rect 940 282 976 297
rect 1034 282 1070 297
rect 1128 282 1164 297
rect 1222 282 1258 297
rect 1316 282 1352 297
rect 1410 282 1446 297
rect 1504 282 1540 297
rect 1598 282 1634 297
rect 1796 282 1832 297
rect 1890 282 1926 297
rect 1984 282 2020 297
rect 2087 282 2123 297
rect 79 261 119 282
rect 173 261 213 282
rect 267 261 307 282
rect 361 261 401 282
rect 22 249 401 261
rect 22 215 38 249
rect 72 215 129 249
rect 163 215 223 249
rect 257 215 317 249
rect 351 215 401 249
rect 22 203 401 215
rect 89 177 119 203
rect 183 177 213 203
rect 277 177 307 203
rect 371 177 401 203
rect 458 261 498 282
rect 552 261 592 282
rect 646 261 686 282
rect 740 261 780 282
rect 938 261 978 282
rect 1032 261 1072 282
rect 1126 261 1166 282
rect 1220 261 1260 282
rect 458 249 780 261
rect 458 215 507 249
rect 541 215 601 249
rect 635 215 696 249
rect 730 215 780 249
rect 458 203 780 215
rect 458 177 488 203
rect 552 177 582 203
rect 646 177 676 203
rect 750 177 780 203
rect 834 249 1260 261
rect 834 215 850 249
rect 884 215 944 249
rect 978 215 1038 249
rect 1072 215 1132 249
rect 1166 215 1260 249
rect 834 203 1260 215
rect 1314 261 1354 282
rect 1408 261 1448 282
rect 1502 261 1542 282
rect 1596 261 1636 282
rect 1314 249 1636 261
rect 1314 215 1364 249
rect 1398 215 1458 249
rect 1492 215 1552 249
rect 1586 215 1636 249
rect 1314 203 1636 215
rect 834 177 864 203
rect 928 177 958 203
rect 1022 177 1052 203
rect 1148 177 1178 203
rect 1314 177 1344 203
rect 1408 177 1438 203
rect 1502 177 1532 203
rect 1606 177 1636 203
rect 1794 261 1834 282
rect 1888 261 1928 282
rect 1982 261 2022 282
rect 2085 261 2125 282
rect 1794 249 2166 261
rect 1794 215 1844 249
rect 1878 215 1938 249
rect 1972 215 2032 249
rect 2066 215 2106 249
rect 2140 215 2166 249
rect 1794 203 2166 215
rect 1794 177 1824 203
rect 1888 177 1918 203
rect 1982 177 2012 203
rect 2085 177 2115 203
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 458 21 488 47
rect 552 21 582 47
rect 646 21 676 47
rect 750 21 780 47
rect 834 21 864 47
rect 928 21 958 47
rect 1022 21 1052 47
rect 1148 21 1178 47
rect 1314 21 1344 47
rect 1408 21 1438 47
rect 1502 21 1532 47
rect 1606 21 1636 47
rect 1794 21 1824 47
rect 1888 21 1918 47
rect 1982 21 2012 47
rect 2085 21 2115 47
<< polycont >>
rect 38 215 72 249
rect 129 215 163 249
rect 223 215 257 249
rect 317 215 351 249
rect 507 215 541 249
rect 601 215 635 249
rect 696 215 730 249
rect 850 215 884 249
rect 944 215 978 249
rect 1038 215 1072 249
rect 1132 215 1166 249
rect 1364 215 1398 249
rect 1458 215 1492 249
rect 1552 215 1586 249
rect 1844 215 1878 249
rect 1938 215 1972 249
rect 2032 215 2066 249
rect 2106 215 2140 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 18 485 448 493
rect 18 451 35 485
rect 69 451 223 485
rect 257 451 448 485
rect 18 417 69 451
rect 223 417 257 451
rect 482 485 558 527
rect 670 485 746 527
rect 482 451 508 485
rect 542 451 558 485
rect 482 435 558 451
rect 602 469 636 485
rect 670 451 696 485
rect 730 451 746 485
rect 670 435 746 451
rect 790 469 840 493
rect 824 435 840 469
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 223 367 257 383
rect 291 383 317 417
rect 351 383 370 417
rect 103 315 129 349
rect 163 333 179 349
rect 291 349 370 383
rect 414 401 448 417
rect 602 401 636 435
rect 790 401 840 435
rect 414 367 602 401
rect 636 367 790 401
rect 824 367 840 401
rect 878 485 1696 493
rect 878 451 894 485
rect 928 451 1082 485
rect 1116 451 1270 485
rect 1304 451 1458 485
rect 1492 451 1646 485
rect 1680 451 1696 485
rect 878 417 928 451
rect 1082 417 1116 451
rect 1270 417 1304 451
rect 1458 417 1492 451
rect 1646 417 1696 451
rect 878 383 894 417
rect 878 367 928 383
rect 972 383 988 417
rect 1022 383 1038 417
rect 291 333 317 349
rect 163 315 317 333
rect 351 333 370 349
rect 972 349 1038 383
rect 1082 367 1116 383
rect 1150 383 1176 417
rect 1210 383 1226 417
rect 972 333 988 349
rect 351 315 988 333
rect 1022 333 1038 349
rect 1150 349 1226 383
rect 1270 367 1304 383
rect 1338 383 1364 417
rect 1398 383 1414 417
rect 1150 333 1176 349
rect 1022 315 1176 333
rect 1210 315 1226 349
rect 103 299 1226 315
rect 1338 349 1414 383
rect 1458 367 1492 383
rect 1526 383 1552 417
rect 1586 383 1602 417
rect 1338 315 1364 349
rect 1398 333 1414 349
rect 1526 349 1602 383
rect 1680 383 1696 417
rect 1646 367 1696 383
rect 1734 485 1784 527
rect 1734 451 1750 485
rect 1734 417 1784 451
rect 1734 383 1750 417
rect 1734 367 1784 383
rect 1818 485 1894 493
rect 1818 451 1844 485
rect 1878 451 1894 485
rect 1818 417 1894 451
rect 1818 383 1844 417
rect 1878 383 1894 417
rect 1526 333 1552 349
rect 1398 315 1552 333
rect 1586 333 1602 349
rect 1818 349 1894 383
rect 1938 485 1972 527
rect 1938 417 1972 451
rect 1938 367 1972 383
rect 2006 485 2082 493
rect 2006 451 2032 485
rect 2066 451 2082 485
rect 2006 417 2082 451
rect 2006 383 2032 417
rect 2066 383 2082 417
rect 1818 333 1844 349
rect 1586 315 1844 333
rect 1878 333 1894 349
rect 2006 349 2082 383
rect 2006 333 2032 349
rect 1878 315 2032 333
rect 2066 315 2082 349
rect 1338 299 2082 315
rect 2135 485 2185 527
rect 2169 451 2185 485
rect 2135 417 2185 451
rect 2169 383 2185 417
rect 2135 349 2185 383
rect 2169 315 2185 349
rect 2135 299 2185 315
rect 22 249 367 255
rect 22 215 38 249
rect 72 215 129 249
rect 163 215 223 249
rect 257 215 317 249
rect 351 215 367 249
rect 411 181 447 299
rect 481 249 788 255
rect 481 215 507 249
rect 541 215 601 249
rect 635 215 696 249
rect 730 215 788 249
rect 834 249 1196 255
rect 834 215 850 249
rect 884 215 944 249
rect 978 215 1038 249
rect 1072 215 1132 249
rect 1166 215 1196 249
rect 1304 249 1602 255
rect 1304 215 1364 249
rect 1398 215 1458 249
rect 1492 215 1552 249
rect 1586 215 1602 249
rect 1818 249 2185 255
rect 1818 215 1844 249
rect 1878 215 1938 249
rect 1972 215 2032 249
rect 2066 215 2106 249
rect 2140 215 2185 249
rect 18 161 69 181
rect 18 127 35 161
rect 103 165 746 181
rect 103 131 129 165
rect 163 131 317 165
rect 351 131 508 165
rect 542 131 696 165
rect 730 131 746 165
rect 790 165 2185 181
rect 824 147 978 165
rect 824 131 840 147
rect 18 93 69 127
rect 790 93 840 131
rect 952 131 978 147
rect 1012 147 1198 165
rect 1012 131 1028 147
rect 18 59 35 93
rect 69 59 223 93
rect 257 59 411 93
rect 445 59 602 93
rect 636 59 790 93
rect 824 59 840 93
rect 18 51 840 59
rect 884 93 918 109
rect 884 17 918 59
rect 952 93 1028 131
rect 1182 131 1198 147
rect 1232 131 1266 165
rect 1300 147 1458 165
rect 1300 131 1316 147
rect 952 59 978 93
rect 1012 59 1028 93
rect 952 51 1028 59
rect 1072 93 1138 109
rect 1072 59 1088 93
rect 1122 59 1138 93
rect 1072 17 1138 59
rect 1182 93 1316 131
rect 1432 131 1458 147
rect 1492 147 1646 165
rect 1492 131 1508 147
rect 1182 59 1198 93
rect 1232 59 1266 93
rect 1300 59 1316 93
rect 1182 51 1316 59
rect 1364 93 1398 109
rect 1364 17 1398 59
rect 1432 93 1508 131
rect 1620 131 1646 147
rect 1680 131 1718 165
rect 1752 147 1938 165
rect 1752 131 1768 147
rect 1432 59 1458 93
rect 1492 59 1508 93
rect 1432 51 1508 59
rect 1552 93 1586 109
rect 1552 17 1586 59
rect 1620 93 1768 131
rect 1912 131 1938 147
rect 1972 147 2135 165
rect 1972 131 1988 147
rect 1620 59 1646 93
rect 1680 59 1718 93
rect 1752 59 1768 93
rect 1620 51 1768 59
rect 1844 93 1878 109
rect 1844 17 1878 59
rect 1912 93 1988 131
rect 2109 131 2135 147
rect 2169 131 2185 165
rect 1912 59 1938 93
rect 1972 59 1988 93
rect 1912 51 1988 59
rect 2032 93 2075 109
rect 2032 59 2041 93
rect 2032 17 2075 59
rect 2109 93 2185 131
rect 2109 59 2135 93
rect 2169 59 2185 93
rect 2109 51 2185 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel locali s 2052 221 2086 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 2144 221 2178 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 1869 221 1903 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 1962 221 1996 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 1408 221 1442 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 1316 221 1350 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 1499 221 1533 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 1037 221 1071 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 948 221 982 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 1135 221 1169 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 250 0 0 0 B1
port 4 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 250 0 0 0 B1
port 4 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 250 0 0 0 B1
port 4 nsew signal input
flabel locali s 307 357 341 391 0 FreeSans 250 0 0 0 Y
port 10 nsew signal output
flabel locali s 216 221 250 255 0 FreeSans 250 0 0 0 B2
port 5 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 B2
port 5 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 B2
port 5 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o32ai_4
<< properties >>
string FIXED_BBOX 0 0 2208 544
string GDS_END 2211484
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 2194514
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
