magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 9 21 725 203
rect 29 -17 63 21
<< scnmos >>
rect 97 47 127 177
rect 183 47 213 177
rect 287 47 317 177
rect 383 47 413 177
rect 581 47 611 177
<< scpmoshvt >>
rect 89 297 125 497
rect 185 297 221 497
rect 279 297 315 497
rect 375 297 411 497
rect 573 297 609 497
<< ndiff >>
rect 35 95 97 177
rect 35 61 43 95
rect 77 61 97 95
rect 35 47 97 61
rect 127 117 183 177
rect 127 83 137 117
rect 171 83 183 117
rect 127 47 183 83
rect 213 95 287 177
rect 213 61 233 95
rect 267 61 287 95
rect 213 47 287 61
rect 317 47 383 177
rect 413 97 581 177
rect 413 63 423 97
rect 457 63 523 97
rect 557 63 581 97
rect 413 47 581 63
rect 611 168 699 177
rect 611 134 651 168
rect 685 134 699 168
rect 611 100 699 134
rect 611 66 651 100
rect 685 66 699 100
rect 611 47 699 66
<< pdiff >>
rect 35 485 89 497
rect 35 451 43 485
rect 77 451 89 485
rect 35 417 89 451
rect 35 383 43 417
rect 77 383 89 417
rect 35 297 89 383
rect 125 297 185 497
rect 221 475 279 497
rect 221 441 233 475
rect 267 441 279 475
rect 221 407 279 441
rect 221 373 233 407
rect 267 373 279 407
rect 221 297 279 373
rect 315 475 375 497
rect 315 441 327 475
rect 361 441 375 475
rect 315 407 375 441
rect 315 373 327 407
rect 361 373 375 407
rect 315 297 375 373
rect 411 475 465 497
rect 411 441 423 475
rect 457 441 465 475
rect 411 297 465 441
rect 519 475 573 497
rect 519 441 527 475
rect 561 441 573 475
rect 519 407 573 441
rect 519 373 527 407
rect 561 373 573 407
rect 519 297 573 373
rect 609 477 699 497
rect 609 443 649 477
rect 683 443 699 477
rect 609 409 699 443
rect 609 375 649 409
rect 683 375 699 409
rect 609 341 699 375
rect 609 307 649 341
rect 683 307 699 341
rect 609 297 699 307
<< ndiffc >>
rect 43 61 77 95
rect 137 83 171 117
rect 233 61 267 95
rect 423 63 457 97
rect 523 63 557 97
rect 651 134 685 168
rect 651 66 685 100
<< pdiffc >>
rect 43 451 77 485
rect 43 383 77 417
rect 233 441 267 475
rect 233 373 267 407
rect 327 441 361 475
rect 327 373 361 407
rect 423 441 457 475
rect 527 441 561 475
rect 527 373 561 407
rect 649 443 683 477
rect 649 375 683 409
rect 649 307 683 341
<< poly >>
rect 89 497 125 523
rect 185 497 221 523
rect 279 497 315 523
rect 375 497 411 523
rect 573 497 609 523
rect 89 282 125 297
rect 185 282 221 297
rect 279 282 315 297
rect 375 282 411 297
rect 573 282 609 297
rect 87 265 127 282
rect 183 265 223 282
rect 277 265 317 282
rect 373 265 413 282
rect 571 265 611 282
rect 87 249 141 265
rect 87 215 97 249
rect 131 215 141 249
rect 87 199 141 215
rect 183 249 317 265
rect 183 215 224 249
rect 258 215 317 249
rect 183 199 317 215
rect 359 249 413 265
rect 359 215 369 249
rect 403 215 413 249
rect 359 199 413 215
rect 505 249 611 265
rect 505 215 515 249
rect 549 215 611 249
rect 505 199 611 215
rect 97 177 127 199
rect 183 177 213 199
rect 287 177 317 199
rect 383 177 413 199
rect 581 177 611 199
rect 97 21 127 47
rect 183 21 213 47
rect 287 21 317 47
rect 383 21 413 47
rect 581 21 611 47
<< polycont >>
rect 97 215 131 249
rect 224 215 258 249
rect 369 215 403 249
rect 515 215 549 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 485 93 493
rect 17 451 43 485
rect 77 451 93 485
rect 17 417 93 451
rect 17 383 43 417
rect 77 383 93 417
rect 17 357 93 383
rect 233 475 267 527
rect 233 407 267 441
rect 233 357 267 373
rect 301 475 377 493
rect 301 441 327 475
rect 361 441 377 475
rect 301 407 377 441
rect 423 475 457 527
rect 423 425 457 441
rect 491 475 571 493
rect 491 441 527 475
rect 561 441 571 475
rect 301 373 327 407
rect 361 391 377 407
rect 491 407 571 441
rect 491 391 527 407
rect 361 373 527 391
rect 561 373 571 407
rect 301 357 571 373
rect 645 477 709 493
rect 645 443 649 477
rect 683 443 709 477
rect 645 409 709 443
rect 645 375 649 409
rect 683 375 709 409
rect 17 165 51 357
rect 645 341 709 375
rect 85 289 378 323
rect 645 307 649 341
rect 683 307 709 341
rect 85 249 155 289
rect 85 215 97 249
rect 131 215 155 249
rect 191 249 300 255
rect 191 215 224 249
rect 258 215 300 249
rect 344 249 378 289
rect 583 273 709 307
rect 503 249 549 265
rect 344 215 369 249
rect 403 215 431 249
rect 503 215 515 249
rect 85 199 155 215
rect 503 165 549 215
rect 17 131 549 165
rect 137 117 171 131
rect 27 61 43 95
rect 77 61 93 95
rect 583 97 617 273
rect 137 67 171 83
rect 27 17 93 61
rect 207 61 233 95
rect 267 61 283 95
rect 376 63 423 97
rect 457 63 523 97
rect 557 63 617 97
rect 651 168 709 184
rect 685 134 709 168
rect 651 100 709 134
rect 685 66 709 100
rect 207 17 283 61
rect 651 17 709 66
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 131 289 165 323 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 663 289 697 323 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 191 215 300 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 xor2_1
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 2820446
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 2814808
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
