magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 821 201
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 175
rect 161 47 191 175
rect 419 47 449 175
rect 491 47 521 175
rect 597 47 627 175
rect 703 47 733 175
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 411 297 447 497
rect 505 297 541 497
rect 599 297 635 497
rect 705 297 741 497
<< ndiff >>
rect 27 161 89 175
rect 27 127 35 161
rect 69 127 89 161
rect 27 93 89 127
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 47 161 175
rect 191 93 419 175
rect 191 59 211 93
rect 245 59 279 93
rect 313 59 419 93
rect 191 47 419 59
rect 449 47 491 175
rect 521 163 597 175
rect 521 129 545 163
rect 579 129 597 163
rect 521 93 597 129
rect 521 59 545 93
rect 579 59 597 93
rect 521 47 597 59
rect 627 47 703 175
rect 733 161 795 175
rect 733 127 743 161
rect 777 127 795 161
rect 733 93 795 127
rect 733 59 743 93
rect 777 59 795 93
rect 733 47 795 59
<< pdiff >>
rect 27 439 81 497
rect 27 405 35 439
rect 69 405 81 439
rect 27 370 81 405
rect 27 336 35 370
rect 69 336 81 370
rect 27 297 81 336
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 297 175 443
rect 211 343 265 497
rect 211 309 223 343
rect 257 309 265 343
rect 211 297 265 309
rect 357 350 411 497
rect 357 316 365 350
rect 399 316 411 350
rect 357 297 411 316
rect 447 477 505 497
rect 447 443 459 477
rect 493 443 505 477
rect 447 297 505 443
rect 541 424 599 497
rect 541 390 553 424
rect 587 390 599 424
rect 541 350 599 390
rect 541 316 553 350
rect 587 316 599 350
rect 541 297 599 316
rect 635 485 705 497
rect 635 451 647 485
rect 681 451 705 485
rect 635 415 705 451
rect 635 381 647 415
rect 681 381 705 415
rect 635 297 705 381
rect 741 424 795 497
rect 741 390 753 424
rect 787 390 795 424
rect 741 350 795 390
rect 741 316 753 350
rect 787 316 795 350
rect 741 297 795 316
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 211 59 245 93
rect 279 59 313 93
rect 545 129 579 163
rect 545 59 579 93
rect 743 127 777 161
rect 743 59 777 93
<< pdiffc >>
rect 35 405 69 439
rect 35 336 69 370
rect 129 443 163 477
rect 223 309 257 343
rect 365 316 399 350
rect 459 443 493 477
rect 553 390 587 424
rect 553 316 587 350
rect 647 451 681 485
rect 647 381 681 415
rect 753 390 787 424
rect 753 316 787 350
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 411 497 447 523
rect 505 497 541 523
rect 599 497 635 523
rect 705 497 741 523
rect 81 282 117 297
rect 175 282 211 297
rect 411 282 447 297
rect 505 282 541 297
rect 599 282 635 297
rect 705 282 741 297
rect 79 266 119 282
rect 173 266 213 282
rect 409 266 449 282
rect 503 266 543 282
rect 597 266 637 282
rect 703 266 743 282
rect 21 250 119 266
rect 21 216 59 250
rect 93 216 119 250
rect 21 200 119 216
rect 89 175 119 200
rect 161 250 225 266
rect 161 216 171 250
rect 205 216 225 250
rect 161 200 225 216
rect 377 250 449 266
rect 377 216 393 250
rect 427 216 449 250
rect 377 200 449 216
rect 161 175 191 200
rect 419 175 449 200
rect 491 250 547 266
rect 491 216 501 250
rect 535 216 547 250
rect 491 200 547 216
rect 597 250 661 266
rect 597 216 607 250
rect 641 216 661 250
rect 597 200 661 216
rect 703 250 767 266
rect 703 216 713 250
rect 747 216 767 250
rect 703 200 767 216
rect 491 175 521 200
rect 597 175 627 200
rect 703 175 733 200
rect 89 21 119 47
rect 161 21 191 47
rect 419 21 449 47
rect 491 21 521 47
rect 597 21 627 47
rect 703 21 733 47
<< polycont >>
rect 59 216 93 250
rect 171 216 205 250
rect 393 216 427 250
rect 501 216 535 250
rect 607 216 641 250
rect 713 216 747 250
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 113 477 493 493
rect 19 439 69 459
rect 19 405 35 439
rect 113 443 129 477
rect 163 459 459 477
rect 163 443 179 459
rect 113 411 179 443
rect 434 443 459 459
rect 631 485 697 527
rect 631 451 647 485
rect 681 451 697 485
rect 434 427 493 443
rect 537 424 587 450
rect 19 370 69 405
rect 19 336 35 370
rect 537 390 553 424
rect 537 366 587 390
rect 631 415 697 451
rect 631 381 647 415
rect 681 381 697 415
rect 753 424 805 450
rect 787 390 805 424
rect 69 343 331 359
rect 69 336 223 343
rect 19 309 223 336
rect 257 309 331 343
rect 19 297 331 309
rect 365 350 587 366
rect 399 316 553 350
rect 753 350 805 390
rect 587 316 753 347
rect 787 316 805 350
rect 365 300 805 316
rect 17 250 119 263
rect 17 216 59 250
rect 93 216 119 250
rect 17 200 119 216
rect 153 250 247 263
rect 153 216 171 250
rect 205 216 247 250
rect 153 200 247 216
rect 281 163 331 297
rect 377 250 449 266
rect 377 216 393 250
rect 427 216 449 250
rect 377 200 449 216
rect 483 250 547 266
rect 483 216 501 250
rect 535 216 547 250
rect 483 200 547 216
rect 581 250 661 266
rect 581 216 607 250
rect 641 216 661 250
rect 581 200 661 216
rect 695 250 799 266
rect 695 216 713 250
rect 747 216 799 250
rect 695 200 799 216
rect 19 161 545 163
rect 19 127 35 161
rect 69 129 545 161
rect 579 129 595 163
rect 69 127 85 129
rect 19 93 85 127
rect 482 93 595 129
rect 19 59 35 93
rect 69 59 85 93
rect 19 51 85 59
rect 185 59 211 93
rect 245 59 279 93
rect 313 59 341 93
rect 482 59 545 93
rect 579 59 595 93
rect 711 161 793 163
rect 711 127 743 161
rect 777 127 793 161
rect 711 93 793 127
rect 711 59 743 93
rect 777 59 793 93
rect 185 17 341 59
rect 711 17 793 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a222oi_1
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 7 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 10 nsew power bidirectional
flabel locali s 174 218 218 252 0 FreeSans 340 0 0 0 C2
port 6 nsew signal input
flabel locali s 31 218 65 252 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 494 218 528 252 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 759 214 793 248 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 587 218 621 252 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 281 218 315 252 0 FreeSans 340 0 0 0 Y
port 11 nsew signal output
flabel locali s 397 218 431 252 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 494 85 528 119 0 FreeSans 340 0 0 0 Y
port 11 nsew signal output
flabel locali s 34 85 68 119 0 FreeSans 340 0 0 0 Y
port 11 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 329626
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 322542
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
