magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 703 203
rect 29 -17 63 21
<< scnmos >>
rect 93 47 123 177
rect 179 47 209 177
rect 285 47 315 177
rect 357 47 387 177
rect 463 47 493 177
rect 557 47 587 177
<< scpmoshvt >>
rect 85 297 121 497
rect 181 297 217 497
rect 277 297 313 497
rect 371 297 407 497
rect 465 297 501 497
rect 559 297 595 497
<< ndiff >>
rect 27 157 93 177
rect 27 123 39 157
rect 73 123 93 157
rect 27 89 93 123
rect 27 55 39 89
rect 73 55 93 89
rect 27 47 93 55
rect 123 47 179 177
rect 209 157 285 177
rect 209 123 230 157
rect 264 123 285 157
rect 209 89 285 123
rect 209 55 230 89
rect 264 55 285 89
rect 209 47 285 55
rect 315 47 357 177
rect 387 89 463 177
rect 387 55 408 89
rect 442 55 463 89
rect 387 47 463 55
rect 493 169 557 177
rect 493 135 513 169
rect 547 135 557 169
rect 493 101 557 135
rect 493 67 513 101
rect 547 67 557 101
rect 493 47 557 67
rect 587 165 677 177
rect 587 131 635 165
rect 669 131 677 165
rect 587 93 677 131
rect 587 59 635 93
rect 669 59 677 93
rect 587 47 677 59
<< pdiff >>
rect 27 477 85 497
rect 27 443 38 477
rect 72 443 85 477
rect 27 409 85 443
rect 27 375 38 409
rect 72 375 85 409
rect 27 297 85 375
rect 121 489 181 497
rect 121 455 134 489
rect 168 455 181 489
rect 121 297 181 455
rect 217 477 277 497
rect 217 443 230 477
rect 264 443 277 477
rect 217 405 277 443
rect 217 371 230 405
rect 264 371 277 405
rect 217 297 277 371
rect 313 489 371 497
rect 313 455 325 489
rect 359 455 371 489
rect 313 297 371 455
rect 407 489 465 497
rect 407 455 419 489
rect 453 455 465 489
rect 407 421 465 455
rect 407 387 419 421
rect 453 387 465 421
rect 407 297 465 387
rect 501 407 559 497
rect 501 373 513 407
rect 547 373 559 407
rect 501 339 559 373
rect 501 305 513 339
rect 547 305 559 339
rect 501 297 559 305
rect 595 477 669 497
rect 595 443 627 477
rect 661 443 669 477
rect 595 409 669 443
rect 595 375 627 409
rect 661 375 669 409
rect 595 297 669 375
<< ndiffc >>
rect 39 123 73 157
rect 39 55 73 89
rect 230 123 264 157
rect 230 55 264 89
rect 408 55 442 89
rect 513 135 547 169
rect 513 67 547 101
rect 635 131 669 165
rect 635 59 669 93
<< pdiffc >>
rect 38 443 72 477
rect 38 375 72 409
rect 134 455 168 489
rect 230 443 264 477
rect 230 371 264 405
rect 325 455 359 489
rect 419 455 453 489
rect 419 387 453 421
rect 513 373 547 407
rect 513 305 547 339
rect 627 443 661 477
rect 627 375 661 409
<< poly >>
rect 85 497 121 523
rect 181 497 217 523
rect 277 497 313 523
rect 371 497 407 523
rect 465 497 501 523
rect 559 497 595 523
rect 85 282 121 297
rect 181 282 217 297
rect 277 282 313 297
rect 371 282 407 297
rect 465 282 501 297
rect 559 282 595 297
rect 83 261 123 282
rect 47 249 123 261
rect 47 215 63 249
rect 97 215 123 249
rect 47 203 123 215
rect 93 177 123 203
rect 179 265 219 282
rect 275 265 315 282
rect 369 265 409 282
rect 179 249 315 265
rect 179 215 189 249
rect 223 215 267 249
rect 301 215 315 249
rect 179 199 315 215
rect 179 177 209 199
rect 285 177 315 199
rect 357 249 421 265
rect 357 215 367 249
rect 401 215 421 249
rect 357 199 421 215
rect 463 261 503 282
rect 557 261 597 282
rect 463 249 657 261
rect 463 215 607 249
rect 641 215 657 249
rect 463 203 657 215
rect 357 177 387 199
rect 463 177 493 203
rect 557 177 587 203
rect 93 21 123 47
rect 179 21 209 47
rect 285 21 315 47
rect 357 21 387 47
rect 463 21 493 47
rect 557 21 587 47
<< polycont >>
rect 63 215 97 249
rect 189 215 223 249
rect 267 215 301 249
rect 367 215 401 249
rect 607 215 641 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 22 477 74 493
rect 22 443 38 477
rect 72 443 74 477
rect 108 489 184 527
rect 108 455 134 489
rect 168 455 184 489
rect 230 477 264 493
rect 22 421 74 443
rect 230 421 264 443
rect 325 489 359 527
rect 325 439 359 455
rect 403 489 678 493
rect 403 455 419 489
rect 453 477 678 489
rect 453 457 627 477
rect 453 455 469 457
rect 22 409 264 421
rect 22 375 38 409
rect 72 405 264 409
rect 403 421 469 455
rect 617 443 627 457
rect 661 443 678 477
rect 403 405 419 421
rect 72 375 230 405
rect 22 371 230 375
rect 264 387 419 405
rect 453 387 469 421
rect 264 371 469 387
rect 503 407 573 423
rect 503 373 513 407
rect 547 373 573 407
rect 503 339 573 373
rect 617 409 678 443
rect 617 375 627 409
rect 661 375 678 409
rect 617 359 678 375
rect 29 299 426 335
rect 29 249 139 299
rect 29 215 63 249
rect 97 215 139 249
rect 29 207 139 215
rect 179 249 315 265
rect 179 215 189 249
rect 223 215 267 249
rect 301 215 315 249
rect 351 249 426 299
rect 503 305 513 339
rect 547 305 573 339
rect 503 266 573 305
rect 351 215 367 249
rect 401 215 426 249
rect 179 199 315 215
rect 20 157 79 173
rect 482 169 573 266
rect 607 249 707 325
rect 641 215 707 249
rect 607 199 707 215
rect 482 157 513 169
rect 20 123 39 157
rect 73 123 79 157
rect 20 89 79 123
rect 20 55 39 89
rect 73 55 79 89
rect 20 17 79 55
rect 201 123 230 157
rect 264 135 513 157
rect 547 135 573 169
rect 264 123 573 135
rect 201 89 280 123
rect 509 101 573 123
rect 201 55 230 89
rect 264 55 280 89
rect 201 51 280 55
rect 382 55 408 89
rect 442 55 458 89
rect 382 17 458 55
rect 509 67 513 101
rect 547 67 573 101
rect 509 51 573 67
rect 619 131 635 165
rect 669 131 685 165
rect 619 93 685 131
rect 619 59 635 93
rect 669 59 685 93
rect 619 17 685 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 616 221 650 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 641 289 675 323 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 76 289 110 323 0 FreeSans 340 180 0 0 A2
port 2 nsew signal input
flabel locali s 179 199 315 265 0 FreeSans 340 180 0 0 A1
port 1 nsew signal input
flabel locali s 539 85 573 119 0 FreeSans 340 180 0 0 Y
port 8 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21oi_2
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 251038
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 244902
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
