magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 2 67 713 203
rect 2 21 483 67
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 187 47 217 177
rect 271 47 301 177
rect 365 47 395 177
rect 595 93 625 177
<< scpmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 597 413 633 497
<< ndiff >>
rect 28 163 83 177
rect 28 129 39 163
rect 73 129 83 163
rect 28 95 83 129
rect 28 61 39 95
rect 73 61 83 95
rect 28 47 83 61
rect 113 163 187 177
rect 113 129 133 163
rect 167 129 187 163
rect 113 95 187 129
rect 113 61 133 95
rect 167 61 187 95
rect 113 47 187 61
rect 217 95 271 177
rect 217 61 227 95
rect 261 61 271 95
rect 217 47 271 61
rect 301 163 365 177
rect 301 129 321 163
rect 355 129 365 163
rect 301 95 365 129
rect 301 61 321 95
rect 355 61 365 95
rect 301 47 365 61
rect 395 163 457 177
rect 395 129 415 163
rect 449 129 457 163
rect 395 95 457 129
rect 395 61 415 95
rect 449 61 457 95
rect 511 153 595 177
rect 511 119 519 153
rect 553 119 595 153
rect 511 93 595 119
rect 625 153 687 177
rect 625 119 645 153
rect 679 119 687 153
rect 625 93 687 119
rect 395 47 457 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 485 179 497
rect 121 451 133 485
rect 167 451 179 485
rect 121 417 179 451
rect 121 383 133 417
rect 167 383 179 417
rect 121 297 179 383
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 409 367 497
rect 309 375 321 409
rect 355 375 367 409
rect 309 341 367 375
rect 309 307 321 341
rect 355 307 367 341
rect 309 297 367 307
rect 403 479 457 497
rect 403 445 415 479
rect 449 445 457 479
rect 403 411 457 445
rect 511 473 597 497
rect 511 439 519 473
rect 553 439 597 473
rect 511 413 597 439
rect 633 479 687 497
rect 633 445 645 479
rect 679 445 687 479
rect 633 413 687 445
rect 403 377 415 411
rect 449 377 457 411
rect 403 343 457 377
rect 403 309 415 343
rect 449 309 457 343
rect 403 297 457 309
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 415 129 449 163
rect 415 61 449 95
rect 519 119 553 153
rect 645 119 679 153
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 451 167 485
rect 133 383 167 417
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 375 355 409
rect 321 307 355 341
rect 415 445 449 479
rect 519 439 553 473
rect 645 445 679 479
rect 415 377 449 411
rect 415 309 449 343
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 597 497 633 523
rect 597 398 633 413
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 83 265 123 282
rect 177 265 217 282
rect 83 249 217 265
rect 83 215 112 249
rect 146 215 217 249
rect 83 199 217 215
rect 83 177 113 199
rect 187 177 217 199
rect 271 265 311 282
rect 365 265 405 282
rect 595 265 635 398
rect 271 249 481 265
rect 271 215 431 249
rect 465 215 481 249
rect 271 199 481 215
rect 595 249 662 265
rect 595 215 608 249
rect 642 215 662 249
rect 595 199 662 215
rect 271 177 301 199
rect 365 177 395 199
rect 595 177 625 199
rect 83 21 113 47
rect 187 21 217 47
rect 271 21 301 47
rect 365 21 395 47
rect 595 21 625 93
<< polycont >>
rect 112 215 146 249
rect 431 215 465 249
rect 608 215 642 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 477 81 493
rect 17 443 39 477
rect 73 443 81 477
rect 17 409 81 443
rect 17 375 39 409
rect 73 375 81 409
rect 17 341 81 375
rect 125 485 175 527
rect 125 451 133 485
rect 167 451 175 485
rect 125 417 175 451
rect 125 383 133 417
rect 167 383 175 417
rect 125 365 175 383
rect 219 479 465 493
rect 219 477 415 479
rect 219 443 227 477
rect 261 459 415 477
rect 261 443 269 459
rect 219 409 269 443
rect 407 445 415 459
rect 449 445 465 479
rect 219 375 227 409
rect 261 375 269 409
rect 17 307 39 341
rect 73 331 81 341
rect 219 341 269 375
rect 219 331 227 341
rect 73 307 227 331
rect 261 307 269 341
rect 17 289 269 307
rect 313 409 363 425
rect 313 375 321 409
rect 355 375 363 409
rect 313 341 363 375
rect 313 307 321 341
rect 355 307 363 341
rect 96 249 252 255
rect 96 215 112 249
rect 146 215 252 249
rect 96 213 252 215
rect 313 179 363 307
rect 407 411 465 445
rect 407 377 415 411
rect 449 377 465 411
rect 407 343 465 377
rect 407 309 415 343
rect 449 309 465 343
rect 407 289 465 309
rect 519 473 553 492
rect 519 249 553 439
rect 637 479 687 527
rect 637 445 645 479
rect 679 445 687 479
rect 637 429 687 445
rect 654 255 707 393
rect 415 215 431 249
rect 465 215 553 249
rect 17 163 73 179
rect 17 129 39 163
rect 17 95 73 129
rect 17 61 39 95
rect 17 17 73 61
rect 107 163 371 179
rect 107 129 133 163
rect 167 145 321 163
rect 167 129 187 145
rect 107 95 187 129
rect 295 129 321 145
rect 355 129 371 163
rect 107 61 133 95
rect 167 61 187 95
rect 107 51 187 61
rect 227 95 261 111
rect 227 17 261 61
rect 295 95 371 129
rect 295 61 321 95
rect 355 61 371 95
rect 295 51 371 61
rect 415 163 449 179
rect 415 95 449 129
rect 519 153 553 215
rect 592 249 707 255
rect 592 215 608 249
rect 642 215 707 249
rect 592 213 707 215
rect 519 89 553 119
rect 637 153 688 169
rect 637 119 645 153
rect 679 119 688 153
rect 415 17 449 61
rect 637 17 688 119
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 654 255 707 393 0 FreeSans 400 0 0 0 B_N
port 2 nsew signal input
flabel locali s 132 221 166 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 306 85 340 119 0 FreeSans 400 0 0 0 Y
port 7 nsew signal output
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor2b_2
rlabel locali s 592 213 707 255 1 B_N
port 2 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 1709332
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1703162
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
