magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 67 1164 203
rect 1 21 966 67
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 183 47 213 177
rect 267 47 297 177
rect 371 47 401 177
rect 566 47 596 177
rect 670 47 700 177
rect 754 47 784 177
rect 848 47 878 177
rect 1046 93 1076 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 568 297 604 497
rect 662 297 698 497
rect 756 297 792 497
rect 850 297 886 497
rect 1048 413 1084 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 183 177
rect 109 129 129 163
rect 163 129 183 163
rect 109 95 183 129
rect 109 61 129 95
rect 163 61 183 95
rect 109 47 183 61
rect 213 95 267 177
rect 213 61 223 95
rect 257 61 267 95
rect 213 47 267 61
rect 297 163 371 177
rect 297 129 317 163
rect 351 129 371 163
rect 297 95 371 129
rect 297 61 317 95
rect 351 61 371 95
rect 297 47 371 61
rect 401 95 453 177
rect 401 61 411 95
rect 445 61 453 95
rect 401 47 453 61
rect 514 95 566 177
rect 514 61 522 95
rect 556 61 566 95
rect 514 47 566 61
rect 596 163 670 177
rect 596 129 616 163
rect 650 129 670 163
rect 596 95 670 129
rect 596 61 616 95
rect 650 61 670 95
rect 596 47 670 61
rect 700 95 754 177
rect 700 61 710 95
rect 744 61 754 95
rect 700 47 754 61
rect 784 163 848 177
rect 784 129 804 163
rect 838 129 848 163
rect 784 95 848 129
rect 784 61 804 95
rect 838 61 848 95
rect 784 47 848 61
rect 878 163 940 177
rect 878 129 898 163
rect 932 129 940 163
rect 878 95 940 129
rect 878 61 898 95
rect 932 61 940 95
rect 994 149 1046 177
rect 994 115 1002 149
rect 1036 115 1046 149
rect 994 93 1046 115
rect 1076 149 1138 177
rect 1076 115 1096 149
rect 1130 115 1138 149
rect 1076 93 1138 115
rect 878 47 940 61
<< pdiff >>
rect 27 479 81 497
rect 27 445 35 479
rect 69 445 81 479
rect 27 411 81 445
rect 27 377 35 411
rect 69 377 81 411
rect 27 343 81 377
rect 27 309 35 343
rect 69 309 81 343
rect 27 297 81 309
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 297 175 375
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 409 269 443
rect 211 375 223 409
rect 257 375 269 409
rect 211 341 269 375
rect 211 307 223 341
rect 257 307 269 341
rect 211 297 269 307
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 409 363 443
rect 305 375 317 409
rect 351 375 363 409
rect 305 297 363 375
rect 399 411 453 497
rect 399 377 411 411
rect 445 377 453 411
rect 399 343 453 377
rect 399 309 411 343
rect 445 309 453 343
rect 399 297 453 309
rect 514 411 568 497
rect 514 377 522 411
rect 556 377 568 411
rect 514 343 568 377
rect 514 309 522 343
rect 556 309 568 343
rect 514 297 568 309
rect 604 477 662 497
rect 604 443 616 477
rect 650 443 662 477
rect 604 409 662 443
rect 604 375 616 409
rect 650 375 662 409
rect 604 297 662 375
rect 698 477 756 497
rect 698 443 710 477
rect 744 443 756 477
rect 698 409 756 443
rect 698 375 710 409
rect 744 375 756 409
rect 698 341 756 375
rect 698 307 710 341
rect 744 307 756 341
rect 698 297 756 307
rect 792 409 850 497
rect 792 375 804 409
rect 838 375 850 409
rect 792 341 850 375
rect 792 307 804 341
rect 838 307 850 341
rect 792 297 850 307
rect 886 477 940 497
rect 886 443 898 477
rect 932 443 940 477
rect 886 409 940 443
rect 994 474 1048 497
rect 994 440 1002 474
rect 1036 440 1048 474
rect 994 413 1048 440
rect 1084 477 1138 497
rect 1084 443 1096 477
rect 1130 443 1138 477
rect 1084 413 1138 443
rect 886 375 898 409
rect 932 375 940 409
rect 886 297 940 375
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 129 129 163 163
rect 129 61 163 95
rect 223 61 257 95
rect 317 129 351 163
rect 317 61 351 95
rect 411 61 445 95
rect 522 61 556 95
rect 616 129 650 163
rect 616 61 650 95
rect 710 61 744 95
rect 804 129 838 163
rect 804 61 838 95
rect 898 129 932 163
rect 898 61 932 95
rect 1002 115 1036 149
rect 1096 115 1130 149
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 129 443 163 477
rect 129 375 163 409
rect 223 443 257 477
rect 223 375 257 409
rect 223 307 257 341
rect 317 443 351 477
rect 317 375 351 409
rect 411 377 445 411
rect 411 309 445 343
rect 522 377 556 411
rect 522 309 556 343
rect 616 443 650 477
rect 616 375 650 409
rect 710 443 744 477
rect 710 375 744 409
rect 710 307 744 341
rect 804 375 838 409
rect 804 307 838 341
rect 898 443 932 477
rect 1002 440 1036 474
rect 1096 443 1130 477
rect 898 375 932 409
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 568 497 604 523
rect 662 497 698 523
rect 756 497 792 523
rect 850 497 886 523
rect 1048 497 1084 523
rect 1048 398 1084 413
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 568 282 604 297
rect 662 282 698 297
rect 756 282 792 297
rect 850 282 886 297
rect 79 265 119 282
rect 173 265 213 282
rect 79 249 213 265
rect 79 215 108 249
rect 142 215 213 249
rect 79 199 213 215
rect 79 177 109 199
rect 183 177 213 199
rect 267 265 307 282
rect 361 265 401 282
rect 267 249 401 265
rect 267 215 330 249
rect 364 215 401 249
rect 267 199 401 215
rect 267 177 297 199
rect 371 177 401 199
rect 566 265 606 282
rect 660 265 700 282
rect 566 249 700 265
rect 566 215 629 249
rect 663 215 700 249
rect 566 199 700 215
rect 566 177 596 199
rect 670 177 700 199
rect 754 265 794 282
rect 848 265 888 282
rect 1046 265 1086 398
rect 754 249 1004 265
rect 754 215 960 249
rect 994 215 1004 249
rect 754 199 1004 215
rect 1046 249 1111 265
rect 1046 215 1057 249
rect 1091 215 1111 249
rect 1046 199 1111 215
rect 754 177 784 199
rect 848 177 878 199
rect 1046 177 1076 199
rect 1046 67 1076 93
rect 79 21 109 47
rect 183 21 213 47
rect 267 21 297 47
rect 371 21 401 47
rect 566 21 596 47
rect 670 21 700 47
rect 754 21 784 47
rect 848 21 878 47
<< polycont >>
rect 108 215 142 249
rect 330 215 364 249
rect 629 215 663 249
rect 960 215 994 249
rect 1057 215 1091 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 479 85 493
rect 17 445 35 479
rect 69 445 85 479
rect 17 411 85 445
rect 17 377 35 411
rect 69 377 85 411
rect 17 343 85 377
rect 129 477 171 527
rect 163 443 171 477
rect 129 409 171 443
rect 163 375 171 409
rect 129 359 171 375
rect 215 477 265 493
rect 215 443 223 477
rect 257 443 265 477
rect 215 409 265 443
rect 215 375 223 409
rect 257 375 265 409
rect 17 309 35 343
rect 69 325 85 343
rect 215 341 265 375
rect 309 477 658 493
rect 309 443 317 477
rect 351 459 616 477
rect 309 409 351 443
rect 650 443 658 477
rect 309 375 317 409
rect 309 359 351 375
rect 385 411 461 425
rect 385 377 411 411
rect 445 377 461 411
rect 215 325 223 341
rect 69 309 223 325
rect 17 307 223 309
rect 257 325 265 341
rect 385 343 461 377
rect 385 325 411 343
rect 257 309 411 325
rect 445 309 461 343
rect 257 307 461 309
rect 17 291 461 307
rect 495 411 572 425
rect 495 377 522 411
rect 556 377 572 411
rect 495 343 572 377
rect 616 409 658 443
rect 650 375 658 409
rect 616 359 658 375
rect 702 477 939 493
rect 702 443 710 477
rect 744 459 898 477
rect 744 443 752 459
rect 702 409 752 443
rect 890 443 898 459
rect 932 443 939 477
rect 702 375 710 409
rect 744 375 752 409
rect 495 309 522 343
rect 556 325 572 343
rect 702 341 752 375
rect 702 325 710 341
rect 556 309 710 325
rect 495 307 710 309
rect 744 307 752 341
rect 495 291 752 307
rect 796 409 846 425
rect 796 375 804 409
rect 838 375 846 409
rect 796 341 846 375
rect 890 409 939 443
rect 890 375 898 409
rect 932 375 939 409
rect 890 359 939 375
rect 973 474 1044 490
rect 973 440 1002 474
rect 1036 440 1044 474
rect 973 407 1044 440
rect 1088 477 1138 527
rect 1088 443 1096 477
rect 1130 443 1138 477
rect 1088 427 1138 443
rect 796 307 804 341
rect 838 325 846 341
rect 838 307 898 325
rect 796 291 898 307
rect 20 249 268 257
rect 20 215 108 249
rect 142 215 268 249
rect 305 249 530 257
rect 305 215 330 249
rect 364 215 530 249
rect 572 249 732 257
rect 572 215 629 249
rect 663 215 732 249
rect 813 215 898 291
rect 973 249 1007 407
rect 1123 257 1177 391
rect 944 215 960 249
rect 994 215 1007 249
rect 1041 249 1177 257
rect 1041 215 1057 249
rect 1091 215 1177 249
rect 813 181 854 215
rect 17 163 69 181
rect 17 129 35 163
rect 17 95 69 129
rect 17 61 35 95
rect 17 17 69 61
rect 103 163 854 181
rect 973 181 1007 215
rect 103 129 129 163
rect 163 145 317 163
rect 163 129 179 145
rect 103 95 179 129
rect 291 129 317 145
rect 351 145 616 163
rect 351 129 367 145
rect 103 61 129 95
rect 163 61 179 95
rect 103 51 179 61
rect 223 95 257 111
rect 223 17 257 61
rect 291 95 367 129
rect 590 129 616 145
rect 650 145 804 163
rect 650 129 666 145
rect 291 61 317 95
rect 351 61 367 95
rect 291 51 367 61
rect 411 95 556 111
rect 445 61 522 95
rect 411 17 556 61
rect 590 95 666 129
rect 778 129 804 145
rect 838 129 854 163
rect 590 61 616 95
rect 650 61 666 95
rect 590 51 666 61
rect 710 95 744 111
rect 710 17 744 61
rect 778 95 854 129
rect 778 61 804 95
rect 838 61 854 95
rect 778 51 854 61
rect 898 163 939 179
rect 932 129 939 163
rect 898 95 939 129
rect 932 61 939 95
rect 973 149 1044 181
rect 973 115 1002 149
rect 1036 115 1044 149
rect 973 76 1044 115
rect 1088 149 1138 165
rect 1088 115 1096 149
rect 1130 115 1138 149
rect 898 17 939 61
rect 1088 17 1138 115
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 1131 221 1165 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 813 215 898 291 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 582 221 616 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 128 221 162 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 309 221 343 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4b_2
rlabel locali s 813 181 854 215 1 Y
port 9 nsew signal output
rlabel locali s 796 325 846 425 1 Y
port 9 nsew signal output
rlabel locali s 796 291 898 325 1 Y
port 9 nsew signal output
rlabel locali s 778 51 854 145 1 Y
port 9 nsew signal output
rlabel locali s 590 51 666 145 1 Y
port 9 nsew signal output
rlabel locali s 291 51 367 145 1 Y
port 9 nsew signal output
rlabel locali s 103 145 854 181 1 Y
port 9 nsew signal output
rlabel locali s 103 51 179 145 1 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 1804962
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1795244
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
