magic
tech sky130A
magscale 1 2
timestamp 1730264365
<< viali >>
rect -1042 1902 -268 1936
rect 806 1902 1580 1936
rect 401 972 435 1006
rect -64 872 -30 906
rect 124 872 158 906
rect 304 872 338 906
rect 492 872 526 906
rect 127 784 161 818
rect 495 772 529 806
rect -1042 216 -686 250
rect 1224 216 1580 250
<< metal1 >>
rect -1174 1936 1712 1972
rect -1174 1902 -1042 1936
rect -268 1902 806 1936
rect 1580 1902 1712 1936
rect -1174 1875 1712 1902
rect -1062 1728 -1052 1794
rect -996 1728 -986 1794
rect -1184 1412 -1174 1478
rect -1118 1412 -1108 1478
rect -1062 1412 -1052 1478
rect -996 1412 -986 1478
rect -955 1466 -905 1740
rect -324 1728 -314 1794
rect -258 1728 -248 1794
rect -314 1656 -258 1728
rect -324 1590 -314 1656
rect -258 1590 -248 1656
rect -1174 424 -1122 1412
rect -407 1322 -355 1425
rect -324 1412 -314 1478
rect -258 1412 -248 1478
rect -417 1270 -407 1322
rect -355 1270 -345 1322
rect -208 1270 -198 1322
rect -146 1270 -136 1322
rect -1052 882 -996 1162
rect -417 1150 -407 1202
rect -355 1150 -345 1202
rect -814 1006 -764 1108
rect -314 1096 -258 1162
rect -198 1006 -146 1270
rect 573 1236 636 1875
rect 786 1728 796 1794
rect 852 1728 862 1794
rect 674 1656 730 1666
rect 674 1590 687 1656
rect 744 1590 754 1656
rect 674 1478 730 1590
rect 664 1412 674 1478
rect 730 1412 740 1478
rect 786 1412 796 1478
rect 852 1412 862 1478
rect 1443 1466 1493 1740
rect 1534 1728 1590 1794
rect 893 1322 945 1424
rect 1524 1412 1534 1478
rect 1590 1412 1600 1478
rect 1646 1412 1656 1478
rect 1712 1412 1722 1478
rect 674 1270 684 1322
rect 736 1270 746 1322
rect 883 1270 893 1322
rect 945 1270 955 1322
rect -82 1184 -72 1236
rect -20 1184 -10 1236
rect 103 1184 113 1236
rect 165 1184 175 1236
rect 379 1184 389 1236
rect 441 1184 451 1236
rect 563 1184 573 1236
rect 625 1184 636 1236
rect 112 1006 447 1012
rect -824 954 -814 1006
rect -758 954 -748 1006
rect -208 954 -198 1006
rect -146 954 -136 1006
rect -1062 830 -1052 882
rect -996 830 -986 882
rect -1052 674 -996 830
rect -814 728 -764 954
rect -91 922 -81 976
rect -14 922 -4 976
rect 112 972 401 1006
rect 435 972 447 1006
rect 112 966 447 972
rect -76 906 -18 922
rect -76 872 -64 906
rect -30 872 -18 906
rect -76 866 -18 872
rect 112 906 170 966
rect 112 872 124 906
rect 158 872 170 906
rect 112 866 170 872
rect 292 906 350 912
rect 292 872 304 906
rect 338 872 350 906
rect 292 824 350 872
rect 456 846 466 912
rect 543 846 553 912
rect 684 882 736 1270
rect 796 1096 852 1162
rect 883 1150 893 1202
rect 945 1150 955 1202
rect 1302 882 1352 1108
rect 1534 1006 1590 1162
rect 1524 954 1534 1006
rect 1590 954 1600 1006
rect 674 830 684 882
rect 736 830 746 882
rect 1286 830 1296 882
rect 1352 830 1362 882
rect 115 818 350 824
rect 115 787 127 818
rect 161 787 350 818
rect 483 806 541 812
rect 483 787 495 806
rect 529 787 541 806
rect -1184 358 -1174 424
rect -1118 358 -1108 424
rect -1072 358 -1062 424
rect -1006 358 -996 424
rect -814 412 -764 686
rect -732 674 -676 740
rect 105 735 115 787
rect 167 778 350 787
rect 167 735 177 778
rect 473 735 483 787
rect 535 735 545 787
rect 1214 674 1270 740
rect 1302 728 1352 830
rect -732 358 -676 424
rect 573 277 636 674
rect 1214 358 1270 424
rect 1302 412 1352 686
rect 1534 674 1590 954
rect 1660 424 1712 1412
rect 1534 358 1544 424
rect 1600 358 1610 424
rect 1646 358 1656 424
rect 1712 358 1722 424
rect -1174 250 1712 277
rect -1174 216 -1042 250
rect -686 216 1224 250
rect 1580 216 1712 250
rect -1174 180 1712 216
<< via1 >>
rect -1052 1728 -996 1794
rect -1174 1412 -1118 1478
rect -1052 1412 -996 1478
rect -314 1728 -258 1794
rect -314 1590 -258 1656
rect -314 1412 -258 1478
rect -407 1270 -355 1322
rect -198 1270 -146 1322
rect -407 1150 -355 1202
rect 796 1728 852 1794
rect 687 1590 744 1656
rect 674 1412 730 1478
rect 796 1412 852 1478
rect 1534 1412 1590 1478
rect 1656 1412 1712 1478
rect 684 1270 736 1322
rect 893 1270 945 1322
rect -72 1184 -20 1236
rect 113 1184 165 1236
rect 389 1184 441 1236
rect 573 1184 625 1236
rect -814 954 -758 1006
rect -198 954 -146 1006
rect -1052 830 -996 882
rect -81 922 -14 976
rect 466 906 543 912
rect 466 872 492 906
rect 492 872 526 906
rect 526 872 543 906
rect 466 846 543 872
rect 893 1150 945 1202
rect 1534 954 1590 1006
rect 684 830 736 882
rect 1296 830 1352 882
rect -1174 358 -1118 424
rect -1062 358 -1006 424
rect 115 784 127 787
rect 127 784 161 787
rect 161 784 167 787
rect 115 735 167 784
rect 483 772 495 787
rect 495 772 529 787
rect 529 772 535 787
rect 483 735 535 772
rect 1544 358 1600 424
rect 1656 358 1712 424
<< metal2 >>
rect -1052 1794 -996 1804
rect -1174 1728 -1052 1794
rect -1052 1718 -996 1728
rect -314 1794 -258 1804
rect -314 1718 -258 1728
rect 796 1794 852 1804
rect 796 1718 852 1728
rect -314 1656 -258 1666
rect 687 1656 744 1666
rect -258 1590 687 1656
rect -314 1580 -258 1590
rect 687 1580 744 1590
rect -1174 1478 -1118 1488
rect -1052 1478 -996 1488
rect -1118 1412 -1052 1478
rect -1174 1402 -1118 1412
rect -1052 1402 -996 1412
rect -314 1478 -258 1488
rect -192 1478 -136 1488
rect -258 1412 -192 1478
rect -314 1402 -258 1412
rect -192 1402 -136 1412
rect 674 1478 730 1488
rect 796 1478 852 1488
rect 730 1412 796 1478
rect 674 1402 730 1412
rect 796 1402 852 1412
rect 1534 1478 1590 1488
rect 1656 1478 1712 1488
rect 1590 1412 1656 1478
rect 1534 1402 1590 1412
rect 1656 1402 1712 1412
rect -407 1322 -355 1332
rect -198 1322 -146 1332
rect -355 1270 -198 1322
rect -407 1260 -355 1270
rect -198 1260 -146 1270
rect 684 1322 736 1332
rect 893 1322 945 1332
rect 736 1270 893 1322
rect 684 1260 736 1270
rect 893 1260 945 1270
rect -72 1236 -20 1246
rect -407 1202 -355 1212
rect -355 1184 -72 1202
rect 113 1236 165 1246
rect -20 1184 113 1202
rect 389 1236 441 1246
rect 165 1184 389 1202
rect 573 1236 625 1246
rect 441 1184 573 1202
rect 893 1202 945 1212
rect 625 1184 893 1202
rect -355 1150 893 1184
rect -407 1140 -355 1150
rect 893 1140 945 1150
rect -814 1006 -758 1016
rect -198 1006 -146 1016
rect 1534 1006 1590 1016
rect -758 954 -198 1006
rect -146 976 1534 1006
rect -146 954 -81 976
rect -814 944 -758 954
rect -198 944 -146 954
rect -14 954 1534 976
rect 1534 944 1590 954
rect -81 912 -14 922
rect 466 912 543 922
rect -1052 882 -996 892
rect -996 846 466 882
rect 684 882 736 892
rect 1296 882 1352 892
rect 543 846 684 882
rect -996 830 684 846
rect 736 830 1296 882
rect -1052 820 -996 830
rect 684 820 736 830
rect 1296 820 1352 830
rect 115 787 167 797
rect -268 735 115 787
rect 115 725 167 735
rect 483 787 535 797
rect 535 735 806 787
rect 483 725 535 735
rect -1174 424 -1118 434
rect -1062 424 -1006 434
rect -1118 358 -1062 424
rect -1174 348 -1118 358
rect -1062 348 -1006 358
rect 1544 424 1600 434
rect 1656 424 1712 434
rect 1600 358 1656 424
rect 1544 348 1600 358
rect 1656 348 1712 358
<< via2 >>
rect 796 1728 852 1794
rect -192 1412 -136 1478
<< metal3 >>
rect 776 1804 872 1815
rect -212 1718 -202 1804
rect -126 1718 -116 1804
rect 776 1718 786 1804
rect 862 1718 872 1804
rect -202 1478 -126 1718
rect 776 1708 872 1718
rect -202 1412 -192 1478
rect -136 1412 -126 1478
rect -202 1407 -126 1412
<< via3 >>
rect -202 1718 -126 1804
rect 786 1794 862 1804
rect 786 1728 796 1794
rect 796 1728 852 1794
rect 852 1728 862 1794
rect 786 1718 862 1728
<< metal4 >>
rect -203 1804 863 1805
rect -203 1718 -202 1804
rect -126 1718 786 1804
rect 862 1718 863 1804
rect -203 1717 863 1718
use sky130_fd_sc_hdll__nand2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hdll/mag
timestamp 1723858470
transform 1 0 -100 0 1 657
box -38 -48 406 592
use sky130_fd_sc_hdll__nand2_1  x2
timestamp 1723858470
transform 1 0 268 0 1 657
box -38 -48 406 592
use sky130_fd_pr__pfet_01v8_R8XU9D  XM1
timestamp 1730240227
transform 0 1 -655 -1 0 1761
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM2
timestamp 1730240227
transform 0 -1 -655 1 0 1445
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM3
timestamp 1730240227
transform 0 1 1193 -1 0 1761
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM4
timestamp 1730240227
transform 0 1 1193 -1 0 1445
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM5
timestamp 1730240227
transform 0 1 -655 -1 0 1129
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_TGNW9T  XM6
timestamp 1730240227
transform 0 -1 -864 1 0 707
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM7
timestamp 1730240227
transform 0 1 -864 -1 0 391
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_R8XU9D  XM8
timestamp 1730240227
transform 0 1 1193 -1 0 1129
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_TGNW9T  XM9
timestamp 1730240227
transform 0 1 1402 -1 0 707
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM10
timestamp 1730240227
transform 0 1 1402 -1 0 391
box -211 -310 211 310
<< labels >>
flabel metal1 -1152 1887 -1096 1953 0 FreeSans 800 0 0 0 VDDA
port 0 nsew
flabel metal1 -1152 193 -1096 259 0 FreeSans 800 0 0 0 VSSA
port 1 nsew
flabel metal2 -1166 1739 -1130 1769 0 FreeSans 800 0 0 0 INN
port 2 nsew
flabel via1 -1166 1429 -1130 1459 0 FreeSans 800 0 0 0 INP
port 3 nsew
flabel metal2 -237 749 -201 779 0 FreeSans 800 0 0 0 OUT
port 4 nsew
flabel metal2 712 749 748 779 0 FreeSans 800 0 0 0 OUTN
port 6 nsew
<< end >>
