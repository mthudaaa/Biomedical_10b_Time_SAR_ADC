magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 859 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 177 47 207 177
rect 271 47 301 177
rect 375 47 405 177
rect 459 47 489 177
rect 553 47 583 177
rect 647 47 677 177
rect 751 47 781 177
<< scpmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 461 297 497 497
rect 555 297 591 497
rect 649 297 685 497
rect 743 297 779 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 177 177
rect 113 129 133 163
rect 167 129 177 163
rect 113 95 177 129
rect 113 61 133 95
rect 167 61 177 95
rect 113 47 177 61
rect 207 95 271 177
rect 207 61 227 95
rect 261 61 271 95
rect 207 47 271 61
rect 301 163 375 177
rect 301 129 321 163
rect 355 129 375 163
rect 301 95 375 129
rect 301 61 321 95
rect 355 61 375 95
rect 301 47 375 61
rect 405 95 459 177
rect 405 61 415 95
rect 449 61 459 95
rect 405 47 459 61
rect 489 163 553 177
rect 489 129 509 163
rect 543 129 553 163
rect 489 95 553 129
rect 489 61 509 95
rect 543 61 553 95
rect 489 47 553 61
rect 583 95 647 177
rect 583 61 603 95
rect 637 61 647 95
rect 583 47 647 61
rect 677 163 751 177
rect 677 129 697 163
rect 731 129 751 163
rect 677 95 751 129
rect 677 61 697 95
rect 731 61 751 95
rect 677 47 751 61
rect 781 95 833 177
rect 781 61 791 95
rect 825 61 833 95
rect 781 47 833 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 485 179 497
rect 121 451 133 485
rect 167 451 179 485
rect 121 417 179 451
rect 121 383 133 417
rect 167 383 179 417
rect 121 297 179 383
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 485 367 497
rect 309 451 321 485
rect 355 451 367 485
rect 309 417 367 451
rect 309 383 321 417
rect 355 383 367 417
rect 309 297 367 383
rect 403 485 461 497
rect 403 451 415 485
rect 449 451 461 485
rect 403 417 461 451
rect 403 383 415 417
rect 449 383 461 417
rect 403 341 461 383
rect 403 307 415 341
rect 449 307 461 341
rect 403 297 461 307
rect 497 409 555 497
rect 497 375 509 409
rect 543 375 555 409
rect 497 341 555 375
rect 497 307 509 341
rect 543 307 555 341
rect 497 297 555 307
rect 591 489 649 497
rect 591 455 603 489
rect 637 455 649 489
rect 591 421 649 455
rect 591 387 603 421
rect 637 387 649 421
rect 591 297 649 387
rect 685 409 743 497
rect 685 375 697 409
rect 731 375 743 409
rect 685 341 743 375
rect 685 307 697 341
rect 731 307 743 341
rect 685 297 743 307
rect 779 485 835 497
rect 779 451 791 485
rect 825 451 835 485
rect 779 417 835 451
rect 779 383 791 417
rect 825 383 835 417
rect 779 297 835 383
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 415 61 449 95
rect 509 129 543 163
rect 509 61 543 95
rect 603 61 637 95
rect 697 129 731 163
rect 697 61 731 95
rect 791 61 825 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 451 167 485
rect 133 383 167 417
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 451 355 485
rect 321 383 355 417
rect 415 451 449 485
rect 415 383 449 417
rect 415 307 449 341
rect 509 375 543 409
rect 509 307 543 341
rect 603 455 637 489
rect 603 387 637 421
rect 697 375 731 409
rect 697 307 731 341
rect 791 451 825 485
rect 791 383 825 417
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 461 497 497 523
rect 555 497 591 523
rect 649 497 685 523
rect 743 497 779 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 461 282 497 297
rect 555 282 591 297
rect 649 282 685 297
rect 743 282 779 297
rect 83 265 123 282
rect 177 265 217 282
rect 271 265 311 282
rect 365 265 405 282
rect 83 249 405 265
rect 83 215 103 249
rect 137 215 181 249
rect 215 215 259 249
rect 293 215 337 249
rect 371 215 405 249
rect 83 199 405 215
rect 83 177 113 199
rect 177 177 207 199
rect 271 177 301 199
rect 375 177 405 199
rect 459 265 499 282
rect 553 265 593 282
rect 647 265 687 282
rect 741 265 781 282
rect 459 249 781 265
rect 459 215 482 249
rect 516 215 560 249
rect 594 215 638 249
rect 672 215 716 249
rect 750 215 781 249
rect 459 199 781 215
rect 459 177 489 199
rect 553 177 583 199
rect 647 177 677 199
rect 751 177 781 199
rect 83 21 113 47
rect 177 21 207 47
rect 271 21 301 47
rect 375 21 405 47
rect 459 21 489 47
rect 553 21 583 47
rect 647 21 677 47
rect 751 21 781 47
<< polycont >>
rect 103 215 137 249
rect 181 215 215 249
rect 259 215 293 249
rect 337 215 371 249
rect 482 215 516 249
rect 560 215 594 249
rect 638 215 672 249
rect 716 215 750 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 477 73 493
rect 18 443 39 477
rect 18 409 73 443
rect 18 375 39 409
rect 18 341 73 375
rect 107 485 183 527
rect 107 451 133 485
rect 167 451 183 485
rect 107 417 183 451
rect 107 383 133 417
rect 167 383 183 417
rect 107 367 183 383
rect 227 477 261 493
rect 227 409 261 443
rect 18 307 39 341
rect 227 341 261 375
rect 295 485 355 527
rect 295 451 321 485
rect 295 417 355 451
rect 295 383 321 417
rect 295 367 355 383
rect 389 489 858 493
rect 389 485 603 489
rect 389 451 415 485
rect 449 459 603 485
rect 449 451 465 459
rect 389 417 465 451
rect 577 455 603 459
rect 637 485 858 489
rect 637 459 791 485
rect 637 455 653 459
rect 389 383 415 417
rect 449 383 465 417
rect 73 307 227 333
rect 389 341 465 383
rect 389 333 415 341
rect 261 307 415 333
rect 449 307 465 341
rect 18 291 465 307
rect 509 409 543 425
rect 577 421 653 455
rect 765 451 791 459
rect 825 451 858 485
rect 577 387 603 421
rect 637 387 653 421
rect 697 409 731 425
rect 509 349 543 375
rect 765 417 858 451
rect 765 383 791 417
rect 825 383 858 417
rect 697 349 731 375
rect 509 341 898 349
rect 543 307 697 341
rect 731 307 898 341
rect 509 289 898 307
rect 28 249 390 255
rect 28 215 103 249
rect 137 215 181 249
rect 215 215 259 249
rect 293 215 337 249
rect 371 215 390 249
rect 464 249 767 255
rect 464 215 482 249
rect 516 215 560 249
rect 594 215 638 249
rect 672 215 716 249
rect 750 215 767 249
rect 819 181 898 289
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 898 181
rect 107 129 133 163
rect 167 145 321 163
rect 167 129 183 145
rect 107 95 183 129
rect 295 129 321 145
rect 355 145 509 163
rect 355 129 371 145
rect 107 61 133 95
rect 167 61 183 95
rect 107 51 183 61
rect 227 95 261 111
rect 227 17 261 61
rect 295 95 371 129
rect 483 129 509 145
rect 543 145 697 163
rect 543 129 559 145
rect 295 61 321 95
rect 355 61 371 95
rect 295 51 371 61
rect 415 95 449 111
rect 415 17 449 61
rect 483 95 559 129
rect 671 129 697 145
rect 731 145 898 163
rect 731 129 747 145
rect 483 61 509 95
rect 543 61 559 95
rect 483 51 559 61
rect 603 95 637 111
rect 603 17 637 61
rect 671 95 747 129
rect 671 61 697 95
rect 731 61 747 95
rect 671 51 747 61
rect 791 95 848 111
rect 825 61 848 95
rect 791 17 848 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 852 289 886 323 0 FreeSans 400 0 0 0 Y
port 7 nsew signal output
flabel locali s 132 221 166 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 642 221 676 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor2_4
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 1686504
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1679042
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
