magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 723 203
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 177
rect 173 47 203 177
rect 381 47 411 177
rect 485 47 515 177
rect 587 47 617 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 373 297 409 497
rect 477 297 513 497
rect 579 297 615 497
<< ndiff >>
rect 27 165 89 177
rect 27 131 35 165
rect 69 131 89 165
rect 27 97 89 131
rect 27 63 35 97
rect 69 63 89 97
rect 27 47 89 63
rect 119 47 173 177
rect 203 93 259 177
rect 203 59 215 93
rect 249 59 259 93
rect 203 47 259 59
rect 313 93 381 177
rect 313 59 321 93
rect 355 59 381 93
rect 313 47 381 59
rect 411 47 485 177
rect 515 89 587 177
rect 515 55 533 89
rect 567 55 587 89
rect 515 47 587 55
rect 617 101 697 177
rect 617 67 655 101
rect 689 67 697 101
rect 617 47 697 67
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 417 175 497
rect 117 383 129 417
rect 163 383 175 417
rect 117 297 175 383
rect 211 343 265 497
rect 211 309 223 343
rect 257 309 265 343
rect 211 297 265 309
rect 319 485 373 497
rect 319 451 327 485
rect 361 451 373 485
rect 319 297 373 451
rect 409 489 477 497
rect 409 455 429 489
rect 463 455 477 489
rect 409 417 477 455
rect 409 383 423 417
rect 457 383 477 417
rect 409 297 477 383
rect 513 489 579 497
rect 513 455 533 489
rect 567 455 579 489
rect 513 421 579 455
rect 513 387 533 421
rect 567 387 579 421
rect 513 297 579 387
rect 615 477 697 497
rect 615 443 655 477
rect 689 443 697 477
rect 615 409 697 443
rect 615 375 655 409
rect 689 375 697 409
rect 615 297 697 375
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 215 59 249 93
rect 321 59 355 93
rect 533 55 567 89
rect 655 67 689 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 383 163 417
rect 223 309 257 343
rect 327 451 361 485
rect 429 455 463 489
rect 423 383 457 417
rect 533 455 567 489
rect 533 387 567 421
rect 655 443 689 477
rect 655 375 689 409
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 373 497 409 523
rect 477 497 513 523
rect 579 497 615 523
rect 81 282 117 297
rect 175 282 211 297
rect 373 282 409 297
rect 477 282 513 297
rect 579 282 615 297
rect 79 265 119 282
rect 65 249 119 265
rect 65 215 75 249
rect 109 215 119 249
rect 65 199 119 215
rect 89 177 119 199
rect 173 265 213 282
rect 371 271 411 282
rect 173 249 227 265
rect 173 215 183 249
rect 217 215 227 249
rect 173 199 227 215
rect 357 249 411 271
rect 475 265 515 282
rect 577 265 617 282
rect 357 215 367 249
rect 401 215 411 249
rect 357 199 411 215
rect 173 177 203 199
rect 381 177 411 199
rect 461 249 515 265
rect 461 215 471 249
rect 505 215 515 249
rect 461 192 515 215
rect 563 249 617 265
rect 563 215 573 249
rect 607 215 617 249
rect 563 199 617 215
rect 485 177 515 192
rect 587 177 617 199
rect 89 21 119 47
rect 173 21 203 47
rect 381 21 411 47
rect 485 21 515 47
rect 587 21 617 47
<< polycont >>
rect 75 215 109 249
rect 183 215 217 249
rect 367 215 401 249
rect 471 215 505 249
rect 573 215 607 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 18 485 85 493
rect 18 451 35 485
rect 69 451 85 485
rect 308 485 379 527
rect 308 451 327 485
rect 361 451 379 485
rect 413 489 479 493
rect 413 455 429 489
rect 463 455 479 489
rect 18 449 85 451
rect 18 417 69 449
rect 413 417 479 455
rect 18 383 35 417
rect 18 349 69 383
rect 113 383 129 417
rect 163 383 423 417
rect 457 383 479 417
rect 517 489 583 527
rect 517 455 533 489
rect 567 455 583 489
rect 517 421 583 455
rect 517 387 533 421
rect 567 387 583 421
rect 655 477 707 493
rect 689 443 707 477
rect 655 409 707 443
rect 113 377 479 383
rect 689 375 707 409
rect 655 357 707 375
rect 18 315 35 349
rect 69 315 223 343
rect 18 309 223 315
rect 257 309 607 343
rect 18 299 607 309
rect 17 249 125 255
rect 17 215 75 249
rect 109 215 125 249
rect 163 249 257 257
rect 163 215 183 249
rect 217 215 257 249
rect 18 165 119 170
rect 18 131 35 165
rect 69 131 119 165
rect 213 135 257 215
rect 305 249 417 257
rect 305 215 367 249
rect 401 215 417 249
rect 305 213 417 215
rect 455 249 525 257
rect 455 215 471 249
rect 505 215 525 249
rect 305 135 349 213
rect 455 196 525 215
rect 573 249 607 299
rect 573 157 607 215
rect 18 97 119 131
rect 18 63 35 97
rect 69 63 119 97
rect 422 123 607 157
rect 422 93 456 123
rect 673 117 707 357
rect 18 17 119 63
rect 174 59 215 93
rect 249 59 321 93
rect 355 59 456 93
rect 655 101 707 117
rect 174 51 456 59
rect 517 55 533 89
rect 567 55 583 89
rect 517 17 583 55
rect 689 67 707 101
rect 655 51 707 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 315 221 349 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 479 221 513 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 661 425 695 459 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 223 221 257 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 315 153 349 187 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 153 257 187 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 661 357 695 391 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a22o_1
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 336176
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 329684
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
