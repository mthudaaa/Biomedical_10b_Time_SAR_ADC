magic
tech sky130A
magscale 1 2
timestamp 1729877160
<< metal3 >>
rect 1394 196 2194 300
rect 880 -4929 1071 -4928
rect 875 -5031 881 -4929
rect 983 -5031 1071 -4929
rect 880 -5032 1071 -5031
rect 1685 -5460 1789 -5272
rect 1457 -5564 2257 -5460
rect 853 -7912 1190 -7808
rect 1685 -7912 1789 -5564
rect 2697 -7912 2801 -5272
rect 853 -13912 957 -7912
rect 1457 -8444 2257 -8340
rect 1457 -9884 2257 -9780
rect 2724 -10072 2977 -9968
rect 1513 -10674 1651 -10478
rect 1857 -10604 2257 -10500
rect 1857 -11220 1961 -10604
rect 1457 -11324 1961 -11220
rect 2139 -11324 2257 -11220
rect 2527 -11369 2617 -11232
rect 2873 -11752 2977 -10072
rect 2702 -11856 2977 -11752
rect 1457 -12045 2257 -11941
rect 1457 -12764 2257 -12660
rect 2697 -13672 2801 -12472
rect 853 -14016 1101 -13912
rect 1457 -14204 2257 -14100
rect 874 -16896 880 -16792
rect 984 -16896 1045 -16792
rect 1457 -17084 2257 -16980
<< via3 >>
rect 881 -5031 983 -4929
rect 880 -16896 984 -16792
<< metal4 >>
rect -13974 746 17499 850
rect -13974 500 -13870 746
rect -12962 504 -12858 746
rect -11950 504 -11846 746
rect -10938 504 -10834 746
rect -9926 504 -9822 746
rect -8914 504 -8810 746
rect -7902 504 -7798 746
rect -6890 504 -6786 746
rect -5878 504 -5774 746
rect -4866 500 -4762 746
rect -3854 504 -3750 746
rect -2842 504 -2738 746
rect -1830 504 -1726 746
rect -818 504 -714 746
rect 194 494 298 746
rect 1205 504 1309 746
rect 2217 504 2321 746
rect 3227 504 3331 746
rect 4239 504 4343 746
rect 5251 504 5355 746
rect 6263 504 6367 746
rect 7275 504 7379 746
rect 8287 504 8391 746
rect 9299 504 9403 746
rect 10311 504 10415 746
rect 11323 504 11427 746
rect 12335 504 12439 746
rect 13347 504 13451 746
rect 14359 504 14463 746
rect 15371 504 15475 746
rect 16383 504 16487 746
rect 17395 504 17499 746
rect 880 -4929 984 -4928
rect 880 -5031 881 -4929
rect 983 -5031 984 -4929
rect 880 -16791 984 -5031
rect 1685 -5032 1789 488
rect 2697 -5032 2801 488
rect 1685 -7912 1789 -5272
rect 2697 -7912 2801 -5272
rect 1685 -9352 1789 -8152
rect 2697 -8700 2801 -8152
rect 2697 -8804 2968 -8700
rect 2697 -9352 2801 -8804
rect 1685 -13672 1789 -12472
rect 2697 -13020 2801 -12472
rect 2864 -13020 2968 -8804
rect 2697 -13124 2968 -13020
rect 2697 -13672 2801 -13124
rect 1685 -16552 1789 -13912
rect 2697 -16552 2801 -13912
rect 879 -16792 985 -16791
rect 879 -16896 880 -16792
rect 984 -16896 985 -16792
rect 879 -16897 985 -16896
rect 1685 -22312 1789 -16792
rect 2697 -22312 2801 -16792
rect -13494 -22492 -13390 -22328
rect -12482 -22492 -12378 -22328
rect -11470 -22492 -11366 -22328
rect -10458 -22492 -10354 -22328
rect -9446 -22492 -9342 -22328
rect -8434 -22492 -8330 -22328
rect -7422 -22492 -7318 -22328
rect -6410 -22492 -6306 -22328
rect -13494 -22596 -6306 -22492
rect -5398 -22492 -5294 -22328
rect -4386 -22492 -4282 -22328
rect -3374 -22492 -3270 -22328
rect -2362 -22492 -2258 -22328
rect -5398 -22596 -2258 -22492
rect -1350 -22492 -1246 -22328
rect -338 -22492 -234 -22328
rect -1350 -22596 -234 -22492
rect 674 -22492 778 -22328
rect 3707 -22492 3811 -22316
rect 674 -22596 3811 -22492
rect 4719 -22492 4823 -22328
rect 5731 -22492 5835 -22328
rect 4719 -22596 5835 -22492
rect 6743 -22492 6847 -22328
rect 9779 -22492 9883 -22328
rect 6743 -22596 9883 -22492
rect 10791 -22492 10895 -22328
rect 11803 -22492 11907 -22328
rect 12815 -22492 12919 -22328
rect 13827 -22492 13931 -22328
rect 14839 -22492 14943 -22328
rect 15851 -22492 15955 -22328
rect 16863 -22492 16967 -22328
rect 17875 -22492 17979 -22310
rect 10791 -22596 17979 -22492
rect -9952 -22984 -9848 -22596
rect -3880 -22820 -3776 -22596
rect -844 -22656 -740 -22596
rect 5225 -22656 5329 -22596
rect -844 -22760 5329 -22656
rect 8261 -22820 8365 -22596
rect -3880 -22924 8365 -22820
rect 14333 -22984 14437 -22596
rect -9952 -23088 14437 -22984
use sky130_fd_pr__cap_mim_m3_1_DURRY3  sky130_fd_pr__cap_mim_m3_1_DURRY3_0
timestamp 1729812420
transform 1 0 1909 0 1 -10912
box -892 -11520 892 11520
use sky130_fd_pr__cap_mim_m3_1_RV4AQU  sky130_fd_pr__cap_mim_m3_1_RV4AQU_1
timestamp 1729760454
transform 1 0 -6692 0 1 -10912
box -7470 -11520 7470 11520
use sky130_fd_pr__cap_mim_m3_1_RV4AQU  sky130_fd_pr__cap_mim_m3_1_RV4AQU_2
timestamp 1729760454
transform 1 0 10509 0 1 -10912
box -7470 -11520 7470 11520
<< labels >>
flabel metal4 2267 646 2267 648 0 FreeSans 1600 0 0 0 VC
port 0 nsew
flabel metal3 1586 -10576 1586 -10576 0 FreeSans 1600 0 0 0 VCM
port 1 nsew
flabel metal3 2566 -11300 2566 -11300 0 FreeSans 1600 0 0 0 SW[0]
port 2 nsew
flabel metal3 1898 -10980 1898 -10980 0 FreeSans 1600 0 0 0 SW[1]
port 3 nsew
flabel metal3 2824 -10018 2824 -10018 0 FreeSans 1600 0 0 0 SW[2]
port 4 nsew
flabel metal4 2922 -12200 2922 -12200 0 FreeSans 1600 0 0 0 SW[3]
port 5 nsew
flabel metal3 858 -13038 858 -13038 0 FreeSans 1600 0 0 0 SW[4]
port 6 nsew
flabel metal4 904 -6972 904 -6972 0 FreeSans 1600 0 0 0 SW[5]
port 7 nsew
flabel metal4 818 -22570 818 -22570 0 FreeSans 1600 0 0 0 SW[6]
port 8 nsew
flabel metal4 1558 -22728 1558 -22728 0 FreeSans 1600 0 0 0 SW[7]
port 9 nsew
flabel metal4 2694 -22882 2694 -22882 0 FreeSans 1600 0 0 0 SW[8]
port 10 nsew
flabel metal4 4062 -23044 4062 -23044 0 FreeSans 1600 0 0 0 SW[9]
port 11 nsew
<< end >>
