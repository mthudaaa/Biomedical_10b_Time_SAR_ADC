magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1064 157
rect 29 -17 63 21
<< scnmos >>
rect 90 47 120 131
rect 186 47 216 131
rect 272 47 302 131
rect 368 47 398 131
rect 464 47 494 131
rect 560 47 590 131
rect 656 47 686 131
rect 752 47 782 131
rect 848 47 878 131
rect 954 47 984 131
<< scpmoshvt >>
rect 82 297 118 497
rect 178 297 214 497
rect 274 297 310 497
rect 370 297 406 497
rect 466 297 502 497
rect 562 297 598 497
rect 658 297 694 497
rect 754 297 790 497
rect 850 297 886 497
rect 946 297 982 497
<< ndiff >>
rect 27 93 90 131
rect 27 59 35 93
rect 69 59 90 93
rect 27 47 90 59
rect 120 106 186 131
rect 120 72 131 106
rect 165 72 186 106
rect 120 47 186 72
rect 216 106 272 131
rect 216 72 227 106
rect 261 72 272 106
rect 216 47 272 72
rect 302 106 368 131
rect 302 72 323 106
rect 357 72 368 106
rect 302 47 368 72
rect 398 97 464 131
rect 398 63 419 97
rect 453 63 464 97
rect 398 47 464 63
rect 494 106 560 131
rect 494 72 515 106
rect 549 72 560 106
rect 494 47 560 72
rect 590 97 656 131
rect 590 63 611 97
rect 645 63 656 97
rect 590 47 656 63
rect 686 106 752 131
rect 686 72 707 106
rect 741 72 752 106
rect 686 47 752 72
rect 782 97 848 131
rect 782 63 803 97
rect 837 63 848 97
rect 782 47 848 63
rect 878 106 954 131
rect 878 72 899 106
rect 933 72 954 106
rect 878 47 954 72
rect 984 97 1038 131
rect 984 63 996 97
rect 1030 63 1038 97
rect 984 47 1038 63
<< pdiff >>
rect 27 441 82 497
rect 27 407 35 441
rect 69 407 82 441
rect 27 355 82 407
rect 27 321 35 355
rect 69 321 82 355
rect 27 297 82 321
rect 118 441 178 497
rect 118 407 131 441
rect 165 407 178 441
rect 118 355 178 407
rect 118 321 131 355
rect 165 321 178 355
rect 118 297 178 321
rect 214 441 274 497
rect 214 407 227 441
rect 261 407 274 441
rect 214 355 274 407
rect 214 321 227 355
rect 261 321 274 355
rect 214 297 274 321
rect 310 441 370 497
rect 310 407 323 441
rect 357 407 370 441
rect 310 355 370 407
rect 310 321 323 355
rect 357 321 370 355
rect 310 297 370 321
rect 406 461 466 497
rect 406 427 419 461
rect 453 427 466 461
rect 406 297 466 427
rect 502 441 562 497
rect 502 407 515 441
rect 549 407 562 441
rect 502 355 562 407
rect 502 321 515 355
rect 549 321 562 355
rect 502 297 562 321
rect 598 461 658 497
rect 598 427 611 461
rect 645 427 658 461
rect 598 297 658 427
rect 694 441 754 497
rect 694 407 707 441
rect 741 407 754 441
rect 694 355 754 407
rect 694 321 707 355
rect 741 321 754 355
rect 694 297 754 321
rect 790 461 850 497
rect 790 427 803 461
rect 837 427 850 461
rect 790 297 850 427
rect 886 441 946 497
rect 886 407 899 441
rect 933 407 946 441
rect 886 355 946 407
rect 886 321 899 355
rect 933 321 946 355
rect 886 297 946 321
rect 982 461 1037 497
rect 982 427 995 461
rect 1029 427 1037 461
rect 982 297 1037 427
<< ndiffc >>
rect 35 59 69 93
rect 131 72 165 106
rect 227 72 261 106
rect 323 72 357 106
rect 419 63 453 97
rect 515 72 549 106
rect 611 63 645 97
rect 707 72 741 106
rect 803 63 837 97
rect 899 72 933 106
rect 996 63 1030 97
<< pdiffc >>
rect 35 407 69 441
rect 35 321 69 355
rect 131 407 165 441
rect 131 321 165 355
rect 227 407 261 441
rect 227 321 261 355
rect 323 407 357 441
rect 323 321 357 355
rect 419 427 453 461
rect 515 407 549 441
rect 515 321 549 355
rect 611 427 645 461
rect 707 407 741 441
rect 707 321 741 355
rect 803 427 837 461
rect 899 407 933 441
rect 899 321 933 355
rect 995 427 1029 461
<< poly >>
rect 82 497 118 523
rect 178 497 214 523
rect 274 497 310 523
rect 370 497 406 523
rect 466 497 502 523
rect 562 497 598 523
rect 658 497 694 523
rect 754 497 790 523
rect 850 497 886 523
rect 946 497 982 523
rect 82 282 118 297
rect 178 282 214 297
rect 274 282 310 297
rect 370 282 406 297
rect 466 282 502 297
rect 562 282 598 297
rect 658 282 694 297
rect 754 282 790 297
rect 850 282 886 297
rect 946 282 982 297
rect 21 249 216 282
rect 21 215 37 249
rect 71 215 216 249
rect 21 180 216 215
rect 90 131 120 180
rect 186 131 216 180
rect 272 265 312 282
rect 368 265 408 282
rect 464 265 504 282
rect 560 265 600 282
rect 656 265 696 282
rect 752 265 792 282
rect 848 265 888 282
rect 944 265 984 282
rect 272 249 984 265
rect 272 215 322 249
rect 356 215 390 249
rect 424 215 468 249
rect 502 215 546 249
rect 580 215 624 249
rect 658 215 702 249
rect 736 215 984 249
rect 272 190 984 215
rect 272 131 302 190
rect 368 131 398 190
rect 464 131 494 190
rect 560 131 590 190
rect 656 131 686 190
rect 752 131 782 190
rect 848 131 878 190
rect 954 131 984 190
rect 90 21 120 47
rect 186 21 216 47
rect 272 21 302 47
rect 368 21 398 47
rect 464 21 494 47
rect 560 21 590 47
rect 656 21 686 47
rect 752 21 782 47
rect 848 21 878 47
rect 954 21 984 47
<< polycont >>
rect 37 215 71 249
rect 322 215 356 249
rect 390 215 424 249
rect 468 215 502 249
rect 546 215 580 249
rect 624 215 658 249
rect 702 215 736 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 19 441 78 527
rect 19 407 35 441
rect 69 407 78 441
rect 19 355 78 407
rect 19 321 35 355
rect 69 321 78 355
rect 19 305 78 321
rect 124 441 174 492
rect 124 407 131 441
rect 165 407 174 441
rect 124 355 174 407
rect 124 321 131 355
rect 165 321 174 355
rect 124 265 174 321
rect 218 441 270 527
rect 218 407 227 441
rect 261 407 270 441
rect 218 355 270 407
rect 218 321 227 355
rect 261 321 270 355
rect 218 305 270 321
rect 314 441 366 492
rect 314 407 323 441
rect 357 407 366 441
rect 314 355 366 407
rect 410 461 462 527
rect 410 427 419 461
rect 453 427 462 461
rect 410 381 462 427
rect 506 441 558 492
rect 506 407 515 441
rect 549 407 558 441
rect 314 321 323 355
rect 357 347 366 355
rect 506 355 558 407
rect 602 461 654 527
rect 602 427 611 461
rect 645 427 654 461
rect 602 381 654 427
rect 698 441 750 492
rect 698 407 707 441
rect 741 407 750 441
rect 506 347 515 355
rect 357 321 515 347
rect 549 347 558 355
rect 698 355 750 407
rect 794 461 846 527
rect 794 427 803 461
rect 837 427 846 461
rect 794 381 846 427
rect 890 441 942 492
rect 890 407 899 441
rect 933 407 942 441
rect 698 347 707 355
rect 549 321 707 347
rect 741 347 750 355
rect 890 355 942 407
rect 986 461 1045 527
rect 986 427 995 461
rect 1029 427 1045 461
rect 986 381 1045 427
rect 890 347 899 355
rect 741 321 899 347
rect 933 347 942 355
rect 933 321 1046 347
rect 314 299 1046 321
rect 17 249 80 265
rect 17 215 37 249
rect 71 215 80 249
rect 17 143 80 215
rect 124 249 798 265
rect 124 215 322 249
rect 356 215 390 249
rect 424 215 468 249
rect 502 215 546 249
rect 580 215 624 249
rect 658 215 702 249
rect 736 215 798 249
rect 29 93 78 109
rect 29 59 35 93
rect 69 59 78 93
rect 29 17 78 59
rect 124 106 174 215
rect 832 181 1046 299
rect 314 147 1046 181
rect 124 72 131 106
rect 165 72 174 106
rect 124 53 174 72
rect 218 106 270 122
rect 218 72 227 106
rect 261 72 270 106
rect 218 17 270 72
rect 314 106 366 147
rect 314 72 323 106
rect 357 72 366 106
rect 314 56 366 72
rect 410 97 462 113
rect 410 63 419 97
rect 453 63 462 97
rect 410 17 462 63
rect 506 106 558 147
rect 506 72 515 106
rect 549 72 558 106
rect 506 56 558 72
rect 602 97 654 113
rect 602 63 611 97
rect 645 63 654 97
rect 602 17 654 63
rect 698 106 750 147
rect 698 72 707 106
rect 741 72 750 106
rect 698 56 750 72
rect 794 97 846 113
rect 794 63 803 97
rect 837 63 846 97
rect 794 17 846 63
rect 890 106 942 147
rect 890 72 899 106
rect 933 72 942 106
rect 890 56 942 72
rect 986 97 1046 113
rect 986 63 996 97
rect 1030 63 1046 97
rect 986 17 1046 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 949 289 983 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 949 153 983 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 856 153 890 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 856 289 890 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 949 221 983 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 856 221 890 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkbuf_8
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 1055660
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1047454
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
