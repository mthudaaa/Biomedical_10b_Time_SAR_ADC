magic
tech sky130A
magscale 1 2
timestamp 1729978159
<< nwell >>
rect 365 760 528 1081
<< viali >>
rect -1146 1011 -372 1045
rect 523 1011 1297 1045
rect 194 814 228 848
rect -183 710 -116 764
rect -1 714 33 748
rect 110 714 144 748
rect 262 714 329 764
rect 5 626 39 660
rect 230 627 264 661
rect -935 -725 -579 -691
rect 730 -725 1086 -691
<< metal1 >>
rect -1278 1071 -202 1091
rect -1278 1045 -1049 1071
rect -989 1045 -202 1071
rect -1278 1011 -1146 1045
rect -372 1011 -202 1045
rect -1278 995 -202 1011
rect 350 1071 1429 1091
rect 350 1045 1140 1071
rect 1200 1045 1429 1071
rect 350 1011 523 1045
rect 1297 1011 1429 1045
rect 350 995 1429 1011
rect -1278 837 -1222 903
rect -1156 837 -1100 903
rect -519 891 -459 995
rect -1288 663 -1278 729
rect -1222 663 -1212 729
rect -1288 587 -1212 663
rect -1288 521 -1278 587
rect -1222 521 -1212 587
rect -1176 521 -1166 587
rect -1110 521 -1100 587
rect -1059 575 -1009 849
rect -418 837 -362 903
rect -13 848 240 854
rect -13 814 194 848
rect 228 814 240 848
rect -13 808 240 814
rect -310 764 -104 770
rect -310 710 -183 764
rect -116 710 -104 764
rect -310 704 -104 710
rect -13 748 45 808
rect 250 764 461 770
rect -13 714 -1 748
rect 33 714 45 748
rect -13 708 45 714
rect 98 748 156 754
rect 98 714 110 748
rect 144 714 156 748
rect -1288 -518 -1212 521
rect -539 413 -459 533
rect -418 521 -362 587
rect -1059 311 -1049 371
rect -989 311 -979 371
rect -539 353 -529 413
rect -469 353 -459 413
rect -539 343 -459 353
rect -310 413 -230 704
rect 98 666 156 714
rect 250 714 262 764
rect 329 714 461 764
rect 250 708 461 714
rect -7 660 156 666
rect -7 627 5 660
rect 39 627 156 660
rect -17 575 -7 627
rect 45 620 156 627
rect 218 661 276 667
rect 218 627 230 661
rect 264 627 276 661
rect 45 575 55 620
rect 218 575 228 627
rect 280 575 290 627
rect -310 353 -300 413
rect -240 353 -230 413
rect -1059 294 -979 311
rect -310 271 -230 353
rect -1156 205 -1100 271
rect -781 37 -731 211
rect -796 -23 -786 37
rect -726 -23 -716 37
rect -945 -267 -889 -201
rect -781 -207 -731 -23
rect -418 -201 -372 271
rect -310 205 -299 271
rect -243 205 -230 271
rect -310 37 -230 205
rect -310 -23 -300 37
rect -240 -23 -230 37
rect -1288 -584 -1278 -518
rect -1222 -584 -1212 -518
rect -965 -583 -955 -517
rect -899 -583 -889 -517
rect -781 -523 -731 -261
rect -625 -267 -615 -201
rect -559 -267 -549 -201
rect -438 -267 -428 -201
rect -372 -267 -362 -201
rect -418 -277 -372 -267
rect -857 -665 -797 -571
rect -625 -583 -569 -517
rect 45 -665 105 516
rect 381 413 461 708
rect 492 729 568 903
rect 610 891 670 995
rect 492 663 502 729
rect 558 663 568 729
rect 513 521 569 587
rect 1160 575 1210 849
rect 1251 837 1307 903
rect 1364 587 1440 588
rect 381 353 391 413
rect 451 353 461 413
rect 610 413 690 527
rect 1251 521 1261 587
rect 1317 521 1327 587
rect 1363 521 1373 587
rect 1429 521 1440 587
rect 610 353 620 413
rect 680 353 690 413
rect 381 37 461 353
rect 1130 311 1140 371
rect 1200 311 1210 371
rect 1130 280 1210 311
rect 493 205 503 271
rect 559 205 569 271
rect 381 -23 391 37
rect 451 -23 461 37
rect 381 -201 461 -23
rect 523 -201 569 205
rect 883 37 933 211
rect 1251 205 1307 271
rect 868 -23 878 37
rect 938 -23 948 37
rect 381 -267 393 -201
rect 449 -267 461 -201
rect 513 -267 523 -201
rect 579 -267 589 -201
rect 700 -267 710 -201
rect 766 -267 776 -201
rect 883 -207 933 -23
rect 381 -277 461 -267
rect 523 -277 569 -267
rect 720 -583 776 -517
rect 883 -523 933 -261
rect 1040 -267 1096 -201
rect 1364 -517 1440 521
rect 948 -665 1008 -571
rect 1040 -583 1050 -517
rect 1106 -583 1116 -517
rect 1364 -583 1374 -517
rect 1430 -583 1440 -517
rect -1279 -691 1428 -665
rect -1279 -725 -935 -691
rect -579 -725 730 -691
rect 1086 -725 1428 -691
rect -1279 -761 1428 -725
<< via1 >>
rect -1049 1045 -989 1071
rect -1049 1011 -989 1045
rect 1140 1045 1200 1071
rect 1140 1011 1200 1045
rect -1222 837 -1156 903
rect -1278 663 -1222 729
rect -1278 521 -1222 587
rect -1166 521 -1110 587
rect -1049 311 -989 371
rect -529 353 -469 413
rect -7 626 5 627
rect 5 626 39 627
rect 39 626 45 627
rect -7 575 45 626
rect 228 575 280 627
rect -300 353 -240 413
rect -786 -23 -726 37
rect -299 205 -243 271
rect -300 -23 -240 37
rect -1278 -584 -1222 -518
rect -955 -583 -899 -517
rect -615 -267 -559 -201
rect -428 -267 -372 -201
rect 502 663 558 729
rect 391 353 451 413
rect 1261 521 1317 587
rect 1373 521 1429 587
rect 620 353 680 413
rect 1140 311 1200 371
rect 503 205 559 271
rect 391 -23 451 37
rect 878 -23 938 37
rect 393 -267 449 -201
rect 523 -267 579 -201
rect 710 -267 766 -201
rect 1050 -583 1106 -517
rect 1374 -583 1430 -517
<< metal2 >>
rect -1049 1071 -989 1081
rect -1049 1001 -989 1011
rect 1140 1071 1200 1081
rect 1140 1001 1200 1011
rect -1222 903 427 913
rect -1156 837 361 903
rect -1222 827 427 837
rect -1278 729 558 739
rect -1222 666 502 729
rect -1278 653 -1222 663
rect 502 653 558 663
rect -7 627 45 637
rect -1278 587 -1110 597
rect -1222 521 -1166 587
rect -1278 511 -1110 521
rect -539 413 -240 423
rect -1049 371 -989 381
rect -539 353 -529 413
rect -469 353 -300 413
rect -7 405 45 575
rect 228 627 280 637
rect 228 405 280 575
rect 361 587 1429 597
rect 427 521 1261 587
rect 1317 521 1373 587
rect 361 511 1429 521
rect -59 353 45 405
rect 176 353 280 405
rect 391 413 690 423
rect 451 353 620 413
rect 680 353 690 413
rect -539 343 -240 353
rect 391 343 690 353
rect 1140 371 1200 381
rect -1049 301 -989 311
rect 1140 301 1200 311
rect -299 271 559 281
rect -243 205 503 271
rect -299 195 559 205
rect -787 37 -240 47
rect -787 -23 -786 37
rect -726 -23 -300 37
rect -787 -33 -240 -23
rect 391 37 938 47
rect 451 -23 878 37
rect 391 -33 938 -23
rect -615 -201 449 -191
rect -559 -267 -428 -201
rect -372 -267 393 -201
rect -615 -277 449 -267
rect 523 -201 766 -191
rect 579 -267 710 -201
rect 523 -277 766 -267
rect -1278 -517 -899 -507
rect -1278 -518 -955 -517
rect -1222 -583 -955 -518
rect -1222 -584 -899 -583
rect -1278 -594 -899 -584
rect 1050 -517 1430 -507
rect 1106 -583 1374 -517
rect 1050 -593 1430 -583
<< via2 >>
rect -1049 1011 -989 1071
rect 1140 1011 1200 1071
rect 361 837 427 903
rect -1049 311 -989 371
rect 361 521 427 587
rect 1140 311 1200 371
<< metal3 >>
rect -1059 1071 -979 1076
rect -1059 1011 -1049 1071
rect -989 1011 -979 1071
rect -1059 371 -979 1011
rect 1130 1071 1210 1076
rect 1130 1011 1140 1071
rect 1200 1011 1210 1071
rect 351 903 437 908
rect 351 837 361 903
rect 427 837 437 903
rect 351 832 437 837
rect 352 592 437 832
rect 351 587 437 592
rect 351 521 361 587
rect 427 521 437 587
rect 351 516 437 521
rect -1059 311 -1049 371
rect -989 311 -979 371
rect -1059 306 -979 311
rect 1130 371 1210 1011
rect 1130 311 1140 371
rect 1200 311 1210 371
rect 1130 306 1210 311
use sky130_fd_sc_hd__nand2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 -202 0 1 499
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x2
timestamp 1723858470
transform 1 0 74 0 1 499
box -38 -48 314 592
use sky130_fd_pr__pfet_01v8_R8XU9D  XM1
timestamp 1729969613
transform 0 1 -759 -1 0 870
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM2
timestamp 1729969613
transform 0 1 -759 -1 0 554
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM3
timestamp 1729969613
transform 0 1 910 -1 0 870
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM4
timestamp 1729969613
transform 0 1 910 -1 0 554
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM5
timestamp 1729969613
transform 0 1 -759 -1 0 238
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_TGNW9T  XM6
timestamp 1729969613
transform 0 -1 -757 1 0 -234
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM7
timestamp 1729969613
transform 0 -1 -757 1 0 -550
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_R8XU9D  XM8
timestamp 1729969613
transform 0 1 910 -1 0 238
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_TGNW9T  XM9
timestamp 1729969613
transform 0 1 908 -1 0 -234
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM10
timestamp 1729969613
transform 0 1 908 -1 0 -550
box -211 -310 211 310
<< labels >>
flabel metal1 -1256 1017 -1199 1069 0 FreeSans 400 0 0 0 vdda
port 0 nsew
flabel metal1 -1266 845 -1209 897 0 FreeSans 400 0 0 0 inn
port 1 nsew
flabel metal1 -1257 -733 -1200 -681 0 FreeSans 400 0 0 0 vssa
port 3 nsew
flabel metal2 -52 364 -20 393 0 FreeSans 400 0 0 0 out
port 4 nsew
flabel metal2 190 371 222 400 0 FreeSans 400 0 0 0 outn
port 6 nsew
flabel metal1 -1278 379 -1221 431 0 FreeSans 400 0 0 0 inp
port 2 nsew
<< end >>
