magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1185 203
rect 30 -17 64 21
<< scnmos >>
rect 80 47 110 177
rect 176 47 206 177
rect 272 47 302 177
rect 368 47 398 177
rect 577 47 607 177
rect 661 47 691 177
rect 782 47 812 177
rect 874 47 904 177
rect 970 47 1000 177
rect 1066 47 1096 177
<< scpmoshvt >>
rect 156 297 192 497
rect 252 297 288 497
rect 348 297 384 497
rect 444 297 480 497
rect 544 297 580 497
rect 650 297 686 497
rect 790 297 826 497
rect 876 297 912 497
rect 972 297 1008 497
rect 1068 297 1104 497
<< ndiff >>
rect 27 93 80 177
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 161 176 177
rect 110 127 131 161
rect 165 127 176 161
rect 110 47 176 127
rect 206 89 272 177
rect 206 55 227 89
rect 261 55 272 89
rect 206 47 272 55
rect 302 159 368 177
rect 302 125 323 159
rect 357 125 368 159
rect 302 47 368 125
rect 398 93 461 177
rect 398 59 419 93
rect 453 59 461 93
rect 398 47 461 59
rect 525 93 577 177
rect 525 59 533 93
rect 567 59 577 93
rect 525 47 577 59
rect 607 169 661 177
rect 607 135 617 169
rect 651 135 661 169
rect 607 47 661 135
rect 691 157 782 177
rect 691 123 727 157
rect 761 123 782 157
rect 691 89 782 123
rect 691 55 727 89
rect 761 55 782 89
rect 691 47 782 55
rect 812 89 874 177
rect 812 55 827 89
rect 861 55 874 89
rect 812 47 874 55
rect 904 157 970 177
rect 904 123 925 157
rect 959 123 970 157
rect 904 47 970 123
rect 1000 89 1066 177
rect 1000 55 1021 89
rect 1055 55 1066 89
rect 1000 47 1066 55
rect 1096 157 1159 177
rect 1096 123 1117 157
rect 1151 123 1159 157
rect 1096 47 1159 123
<< pdiff >>
rect 91 485 156 497
rect 91 451 99 485
rect 133 451 156 485
rect 91 408 156 451
rect 91 374 99 408
rect 133 374 156 408
rect 91 297 156 374
rect 192 477 252 497
rect 192 443 205 477
rect 239 443 252 477
rect 192 385 252 443
rect 192 351 205 385
rect 239 351 252 385
rect 192 297 252 351
rect 288 485 348 497
rect 288 451 301 485
rect 335 451 348 485
rect 288 408 348 451
rect 288 374 301 408
rect 335 374 348 408
rect 288 297 348 374
rect 384 477 444 497
rect 384 443 397 477
rect 431 443 444 477
rect 384 385 444 443
rect 384 351 397 385
rect 431 351 444 385
rect 384 297 444 351
rect 480 485 544 497
rect 480 451 497 485
rect 531 451 544 485
rect 480 297 544 451
rect 580 477 650 497
rect 580 443 593 477
rect 627 443 650 477
rect 580 409 650 443
rect 580 375 593 409
rect 627 375 650 409
rect 580 297 650 375
rect 686 489 790 497
rect 686 455 719 489
rect 753 455 790 489
rect 686 297 790 455
rect 826 297 876 497
rect 912 489 972 497
rect 912 455 925 489
rect 959 455 972 489
rect 912 421 972 455
rect 912 387 925 421
rect 959 387 972 421
rect 912 297 972 387
rect 1008 297 1068 497
rect 1104 489 1163 497
rect 1104 455 1117 489
rect 1151 455 1163 489
rect 1104 421 1163 455
rect 1104 387 1117 421
rect 1151 387 1163 421
rect 1104 297 1163 387
<< ndiffc >>
rect 35 59 69 93
rect 131 127 165 161
rect 227 55 261 89
rect 323 125 357 159
rect 419 59 453 93
rect 533 59 567 93
rect 617 135 651 169
rect 727 123 761 157
rect 727 55 761 89
rect 827 55 861 89
rect 925 123 959 157
rect 1021 55 1055 89
rect 1117 123 1151 157
<< pdiffc >>
rect 99 451 133 485
rect 99 374 133 408
rect 205 443 239 477
rect 205 351 239 385
rect 301 451 335 485
rect 301 374 335 408
rect 397 443 431 477
rect 397 351 431 385
rect 497 451 531 485
rect 593 443 627 477
rect 593 375 627 409
rect 719 455 753 489
rect 925 455 959 489
rect 925 387 959 421
rect 1117 455 1151 489
rect 1117 387 1151 421
<< poly >>
rect 156 497 192 523
rect 252 497 288 523
rect 348 497 384 523
rect 444 497 480 523
rect 544 497 580 523
rect 650 497 686 523
rect 790 497 826 523
rect 876 497 912 523
rect 972 497 1008 523
rect 1068 497 1104 523
rect 156 282 192 297
rect 252 282 288 297
rect 348 282 384 297
rect 444 282 480 297
rect 544 282 580 297
rect 650 282 686 297
rect 790 282 826 297
rect 876 282 912 297
rect 972 282 1008 297
rect 1068 282 1104 297
rect 154 265 194 282
rect 250 265 290 282
rect 346 265 386 282
rect 442 265 482 282
rect 80 249 482 265
rect 80 215 120 249
rect 154 215 198 249
rect 232 215 266 249
rect 300 215 344 249
rect 378 215 422 249
rect 456 215 482 249
rect 80 199 482 215
rect 542 265 582 282
rect 648 265 688 282
rect 788 265 828 282
rect 542 249 691 265
rect 542 215 563 249
rect 597 215 647 249
rect 681 215 691 249
rect 542 199 691 215
rect 743 249 828 265
rect 743 215 759 249
rect 793 215 828 249
rect 743 199 828 215
rect 874 265 914 282
rect 970 265 1010 282
rect 1066 265 1106 282
rect 874 249 1024 265
rect 874 215 884 249
rect 918 215 970 249
rect 1004 215 1024 249
rect 874 199 1024 215
rect 1066 249 1142 265
rect 1066 215 1082 249
rect 1116 215 1142 249
rect 1066 199 1142 215
rect 80 177 110 199
rect 176 177 206 199
rect 272 177 302 199
rect 368 177 398 199
rect 577 177 607 199
rect 661 177 691 199
rect 782 177 812 199
rect 874 177 904 199
rect 970 177 1000 199
rect 1066 177 1096 199
rect 80 21 110 47
rect 176 21 206 47
rect 272 21 302 47
rect 368 21 398 47
rect 577 21 607 47
rect 661 21 691 47
rect 782 21 812 47
rect 874 21 904 47
rect 970 21 1000 47
rect 1066 21 1096 47
<< polycont >>
rect 120 215 154 249
rect 198 215 232 249
rect 266 215 300 249
rect 344 215 378 249
rect 422 215 456 249
rect 563 215 597 249
rect 647 215 681 249
rect 759 215 793 249
rect 884 215 918 249
rect 970 215 1004 249
rect 1082 215 1116 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 83 485 159 527
rect 83 451 99 485
rect 133 451 159 485
rect 83 408 159 451
rect 83 374 99 408
rect 133 374 159 408
rect 203 477 241 493
rect 203 443 205 477
rect 239 443 241 477
rect 203 385 241 443
rect 203 351 205 385
rect 239 351 241 385
rect 275 485 351 527
rect 275 451 301 485
rect 335 451 351 485
rect 275 408 351 451
rect 275 374 301 408
rect 335 374 351 408
rect 395 477 431 493
rect 395 443 397 477
rect 467 485 547 527
rect 467 451 497 485
rect 531 451 547 485
rect 591 477 639 493
rect 395 385 431 443
rect 591 443 593 477
rect 627 443 639 477
rect 703 489 769 527
rect 1091 489 1173 527
rect 703 455 719 489
rect 753 455 769 489
rect 899 455 925 489
rect 959 455 975 489
rect 591 421 639 443
rect 899 421 975 455
rect 591 417 925 421
rect 203 340 241 351
rect 395 351 397 385
rect 395 340 431 351
rect 18 306 431 340
rect 465 409 925 417
rect 465 375 593 409
rect 627 387 925 409
rect 959 387 975 421
rect 1091 455 1117 489
rect 1151 455 1173 489
rect 1091 421 1173 455
rect 1091 387 1117 421
rect 1151 387 1173 421
rect 627 375 975 387
rect 465 366 639 375
rect 18 161 70 306
rect 465 267 513 366
rect 104 249 513 267
rect 104 215 120 249
rect 154 215 198 249
rect 232 215 266 249
rect 300 215 344 249
rect 378 215 422 249
rect 456 215 513 249
rect 547 249 697 323
rect 547 215 563 249
rect 597 215 647 249
rect 681 215 697 249
rect 752 299 1176 341
rect 752 249 823 299
rect 752 215 759 249
rect 793 215 823 249
rect 104 199 513 215
rect 463 174 513 199
rect 752 198 823 215
rect 884 249 1014 265
rect 918 215 970 249
rect 1004 215 1014 249
rect 884 199 1014 215
rect 1082 249 1176 299
rect 1116 215 1176 249
rect 1082 199 1176 215
rect 463 169 677 174
rect 18 127 131 161
rect 165 159 373 161
rect 165 127 323 159
rect 129 125 323 127
rect 357 125 373 159
rect 463 135 617 169
rect 651 135 677 169
rect 463 131 677 135
rect 129 123 373 125
rect 711 123 727 157
rect 761 123 925 157
rect 959 123 1117 157
rect 1151 123 1167 157
rect 711 97 777 123
rect 517 93 777 97
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 211 55 227 89
rect 261 55 277 89
rect 211 17 277 55
rect 403 59 419 93
rect 453 59 469 93
rect 403 17 469 59
rect 517 59 533 93
rect 567 89 777 93
rect 567 59 727 89
rect 517 55 727 59
rect 761 55 777 89
rect 517 51 777 55
rect 811 55 827 89
rect 861 55 879 89
rect 811 17 879 55
rect 995 55 1021 89
rect 1055 55 1071 89
rect 995 17 1071 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 1132 289 1166 323 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 948 221 982 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 581 289 615 323 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 30 153 64 187 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 o21a_4
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 1917378
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1909038
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
