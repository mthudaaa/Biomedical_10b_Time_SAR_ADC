magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 907 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 168 47 198 177
rect 274 47 304 177
rect 401 47 431 177
rect 507 47 537 177
rect 601 47 631 177
rect 695 47 725 177
rect 799 47 829 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 277 297 313 497
rect 403 297 439 497
rect 509 297 545 497
rect 603 297 639 497
rect 697 297 733 497
rect 791 297 827 497
<< ndiff >>
rect 27 101 89 177
rect 27 67 35 101
rect 69 67 89 101
rect 27 47 89 67
rect 119 47 168 177
rect 198 47 274 177
rect 304 47 401 177
rect 431 94 507 177
rect 431 60 461 94
rect 495 60 507 94
rect 431 47 507 60
rect 537 101 601 177
rect 537 67 557 101
rect 591 67 601 101
rect 537 47 601 67
rect 631 94 695 177
rect 631 60 651 94
rect 685 60 695 94
rect 631 47 695 60
rect 725 101 799 177
rect 725 67 745 101
rect 779 67 799 101
rect 725 47 799 67
rect 829 94 881 177
rect 829 60 839 94
rect 873 60 881 94
rect 829 47 881 60
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 297 81 383
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 297 175 375
rect 211 489 277 497
rect 211 455 227 489
rect 261 455 277 489
rect 211 421 277 455
rect 211 387 227 421
rect 261 387 277 421
rect 211 297 277 387
rect 313 477 403 497
rect 313 443 325 477
rect 359 443 403 477
rect 313 409 403 443
rect 313 375 325 409
rect 359 375 403 409
rect 313 297 403 375
rect 439 489 509 497
rect 439 455 461 489
rect 495 455 509 489
rect 439 421 509 455
rect 439 387 461 421
rect 495 387 509 421
rect 439 297 509 387
rect 545 477 603 497
rect 545 443 557 477
rect 591 443 603 477
rect 545 409 603 443
rect 545 375 557 409
rect 591 375 603 409
rect 545 297 603 375
rect 639 485 697 497
rect 639 451 651 485
rect 685 451 697 485
rect 639 417 697 451
rect 639 383 651 417
rect 685 383 697 417
rect 639 297 697 383
rect 733 477 791 497
rect 733 443 745 477
rect 779 443 791 477
rect 733 409 791 443
rect 733 375 745 409
rect 779 375 791 409
rect 733 297 791 375
rect 827 485 881 497
rect 827 451 839 485
rect 873 451 881 485
rect 827 417 881 451
rect 827 383 839 417
rect 873 383 881 417
rect 827 297 881 383
<< ndiffc >>
rect 35 67 69 101
rect 461 60 495 94
rect 557 67 591 101
rect 651 60 685 94
rect 745 67 779 101
rect 839 60 873 94
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 129 443 163 477
rect 129 375 163 409
rect 227 455 261 489
rect 227 387 261 421
rect 325 443 359 477
rect 325 375 359 409
rect 461 455 495 489
rect 461 387 495 421
rect 557 443 591 477
rect 557 375 591 409
rect 651 451 685 485
rect 651 383 685 417
rect 745 443 779 477
rect 745 375 779 409
rect 839 451 873 485
rect 839 383 873 417
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 277 497 313 523
rect 403 497 439 523
rect 509 497 545 523
rect 603 497 639 523
rect 697 497 733 523
rect 791 497 827 523
rect 81 282 117 297
rect 175 282 211 297
rect 277 282 313 297
rect 403 282 439 297
rect 509 282 545 297
rect 603 282 639 297
rect 697 282 733 297
rect 791 282 827 297
rect 79 265 119 282
rect 22 249 119 265
rect 173 265 213 282
rect 275 265 315 282
rect 401 265 441 282
rect 507 265 547 282
rect 601 265 641 282
rect 695 265 735 282
rect 789 265 829 282
rect 173 261 232 265
rect 22 215 32 249
rect 66 215 119 249
rect 22 199 119 215
rect 89 177 119 199
rect 168 249 232 261
rect 168 215 178 249
rect 212 215 232 249
rect 168 199 232 215
rect 274 249 357 265
rect 274 215 303 249
rect 337 215 357 249
rect 274 199 357 215
rect 401 249 465 265
rect 401 215 411 249
rect 445 215 465 249
rect 168 177 198 199
rect 274 177 304 199
rect 401 193 465 215
rect 507 249 829 265
rect 507 215 581 249
rect 615 215 659 249
rect 693 215 737 249
rect 771 215 829 249
rect 507 199 829 215
rect 401 177 431 193
rect 507 177 537 199
rect 601 177 631 199
rect 695 177 725 199
rect 799 177 829 199
rect 89 21 119 47
rect 168 21 198 47
rect 274 21 304 47
rect 401 21 431 47
rect 507 21 537 47
rect 601 21 631 47
rect 695 21 725 47
rect 799 21 829 47
<< polycont >>
rect 32 215 66 249
rect 178 215 212 249
rect 303 215 337 249
rect 411 215 445 249
rect 581 215 615 249
rect 659 215 693 249
rect 737 215 771 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 21 485 77 527
rect 21 451 35 485
rect 69 451 77 485
rect 21 417 77 451
rect 21 383 35 417
rect 69 383 77 417
rect 21 367 77 383
rect 121 477 163 493
rect 121 443 129 477
rect 121 409 163 443
rect 121 375 129 409
rect 211 489 277 527
rect 211 455 227 489
rect 261 455 277 489
rect 211 421 277 455
rect 211 387 227 421
rect 261 387 277 421
rect 321 477 359 493
rect 321 443 325 477
rect 321 409 359 443
rect 121 333 163 375
rect 321 375 325 409
rect 321 333 359 375
rect 445 489 511 527
rect 445 455 461 489
rect 495 455 511 489
rect 445 421 511 455
rect 445 387 461 421
rect 495 387 511 421
rect 445 371 511 387
rect 557 477 607 493
rect 591 443 607 477
rect 557 409 607 443
rect 591 375 607 409
rect 25 249 66 331
rect 25 215 32 249
rect 25 153 66 215
rect 100 299 523 333
rect 100 117 144 299
rect 35 101 144 117
rect 69 67 144 101
rect 178 249 269 265
rect 212 215 269 249
rect 178 84 269 215
rect 303 249 356 265
rect 337 215 356 249
rect 303 85 356 215
rect 397 249 455 265
rect 397 215 411 249
rect 445 215 455 249
rect 489 261 523 299
rect 557 331 607 375
rect 651 485 701 527
rect 685 451 701 485
rect 651 417 701 451
rect 685 383 701 417
rect 651 367 701 383
rect 745 477 779 493
rect 745 409 779 443
rect 813 485 889 527
rect 813 451 839 485
rect 873 451 889 485
rect 813 417 889 451
rect 813 383 839 417
rect 873 383 889 417
rect 745 349 779 375
rect 745 331 891 349
rect 557 297 891 331
rect 489 249 787 261
rect 489 215 581 249
rect 615 215 659 249
rect 693 215 737 249
rect 771 215 787 249
rect 397 146 455 215
rect 840 162 891 297
rect 557 128 891 162
rect 445 94 507 110
rect 35 51 144 67
rect 445 60 461 94
rect 495 60 507 94
rect 445 17 507 60
rect 557 101 591 128
rect 745 101 779 128
rect 557 51 591 67
rect 625 60 651 94
rect 685 60 701 94
rect 625 17 701 60
rect 745 51 779 67
rect 813 60 839 94
rect 873 60 889 94
rect 813 17 889 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 857 153 891 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 857 221 891 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 305 85 339 119 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 213 85 247 119 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 397 153 431 187 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 857 289 891 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 305 153 339 187 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 213 153 247 187 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4_4
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 849922
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 841902
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
