magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 5190 582
<< pwell >>
rect 1 196 469 203
rect 2107 196 3045 203
rect 4683 196 5151 203
rect 1 157 909 196
rect 1667 157 3485 196
rect 4243 157 5151 196
rect 1 40 5151 157
rect 1 21 469 40
rect 982 21 1594 40
rect 2107 21 3045 40
rect 3558 21 4170 40
rect 4683 21 5151 40
rect 29 -17 63 21
rect 2513 -17 2639 21
rect 5089 -17 5123 21
<< scnmos >>
rect 89 47 119 177
rect 173 47 203 177
rect 277 47 307 177
rect 361 47 391 177
rect 549 66 579 170
rect 633 66 663 170
rect 717 66 747 170
rect 801 66 831 170
rect 1060 47 1090 131
rect 1144 47 1174 131
rect 1402 47 1432 131
rect 1486 47 1516 131
rect 1745 66 1775 170
rect 1829 66 1859 170
rect 1913 66 1943 170
rect 1997 66 2027 170
rect 2185 47 2215 177
rect 2269 47 2299 177
rect 2373 47 2403 177
rect 2457 47 2487 177
rect 2665 47 2695 177
rect 2749 47 2779 177
rect 2853 47 2883 177
rect 2937 47 2967 177
rect 3125 66 3155 170
rect 3209 66 3239 170
rect 3293 66 3323 170
rect 3377 66 3407 170
rect 3636 47 3666 131
rect 3720 47 3750 131
rect 3978 47 4008 131
rect 4062 47 4092 131
rect 4321 66 4351 170
rect 4405 66 4435 170
rect 4489 66 4519 170
rect 4573 66 4603 170
rect 4761 47 4791 177
rect 4845 47 4875 177
rect 4949 47 4979 177
rect 5033 47 5063 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 561 311 597 475
rect 655 311 691 475
rect 749 311 785 475
rect 843 311 879 475
rect 1052 325 1088 489
rect 1146 325 1182 489
rect 1394 325 1430 489
rect 1488 325 1524 489
rect 1697 311 1733 475
rect 1791 311 1827 475
rect 1885 311 1921 475
rect 1979 311 2015 475
rect 2177 297 2213 497
rect 2271 297 2307 497
rect 2365 297 2401 497
rect 2459 297 2495 497
rect 2657 297 2693 497
rect 2751 297 2787 497
rect 2845 297 2881 497
rect 2939 297 2975 497
rect 3137 311 3173 475
rect 3231 311 3267 475
rect 3325 311 3361 475
rect 3419 311 3455 475
rect 3628 325 3664 489
rect 3722 325 3758 489
rect 3970 325 4006 489
rect 4064 325 4100 489
rect 4273 311 4309 475
rect 4367 311 4403 475
rect 4461 311 4497 475
rect 4555 311 4591 475
rect 4753 297 4789 497
rect 4847 297 4883 497
rect 4941 297 4977 497
rect 5035 297 5071 497
<< ndiff >>
rect 27 161 89 177
rect 27 127 45 161
rect 79 127 89 161
rect 27 93 89 127
rect 27 59 45 93
rect 79 59 89 93
rect 27 47 89 59
rect 119 161 173 177
rect 119 127 129 161
rect 163 127 173 161
rect 119 93 173 127
rect 119 59 129 93
rect 163 59 173 93
rect 119 47 173 59
rect 203 93 277 177
rect 203 59 223 93
rect 257 59 277 93
rect 203 47 277 59
rect 307 161 361 177
rect 307 127 317 161
rect 351 127 361 161
rect 307 93 361 127
rect 307 59 317 93
rect 351 59 361 93
rect 307 47 361 59
rect 391 93 443 177
rect 391 59 401 93
rect 435 59 443 93
rect 497 135 549 170
rect 497 101 505 135
rect 539 101 549 135
rect 497 66 549 101
rect 579 153 633 170
rect 579 119 589 153
rect 623 119 633 153
rect 579 66 633 119
rect 663 135 717 170
rect 663 101 673 135
rect 707 101 717 135
rect 663 66 717 101
rect 747 153 801 170
rect 747 119 757 153
rect 791 119 801 153
rect 747 66 801 119
rect 831 135 883 170
rect 831 101 841 135
rect 875 101 883 135
rect 831 66 883 101
rect 391 47 443 59
rect 1008 106 1060 131
rect 1008 72 1016 106
rect 1050 72 1060 106
rect 1008 47 1060 72
rect 1090 106 1144 131
rect 1090 72 1100 106
rect 1134 72 1144 106
rect 1090 47 1144 72
rect 1174 106 1226 131
rect 1174 72 1184 106
rect 1218 72 1226 106
rect 1174 47 1226 72
rect 1350 106 1402 131
rect 1350 72 1358 106
rect 1392 72 1402 106
rect 1350 47 1402 72
rect 1432 106 1486 131
rect 1432 72 1442 106
rect 1476 72 1486 106
rect 1432 47 1486 72
rect 1516 106 1568 131
rect 1516 72 1526 106
rect 1560 72 1568 106
rect 1516 47 1568 72
rect 1693 135 1745 170
rect 1693 101 1701 135
rect 1735 101 1745 135
rect 1693 66 1745 101
rect 1775 153 1829 170
rect 1775 119 1785 153
rect 1819 119 1829 153
rect 1775 66 1829 119
rect 1859 135 1913 170
rect 1859 101 1869 135
rect 1903 101 1913 135
rect 1859 66 1913 101
rect 1943 153 1997 170
rect 1943 119 1953 153
rect 1987 119 1997 153
rect 1943 66 1997 119
rect 2027 135 2079 170
rect 2027 101 2037 135
rect 2071 101 2079 135
rect 2027 66 2079 101
rect 2133 93 2185 177
rect 2133 59 2141 93
rect 2175 59 2185 93
rect 2133 47 2185 59
rect 2215 161 2269 177
rect 2215 127 2225 161
rect 2259 127 2269 161
rect 2215 93 2269 127
rect 2215 59 2225 93
rect 2259 59 2269 93
rect 2215 47 2269 59
rect 2299 93 2373 177
rect 2299 59 2319 93
rect 2353 59 2373 93
rect 2299 47 2373 59
rect 2403 161 2457 177
rect 2403 127 2413 161
rect 2447 127 2457 161
rect 2403 93 2457 127
rect 2403 59 2413 93
rect 2447 59 2457 93
rect 2403 47 2457 59
rect 2487 161 2549 177
rect 2487 127 2497 161
rect 2531 127 2549 161
rect 2487 93 2549 127
rect 2487 59 2497 93
rect 2531 59 2549 93
rect 2487 47 2549 59
rect 2603 161 2665 177
rect 2603 127 2621 161
rect 2655 127 2665 161
rect 2603 93 2665 127
rect 2603 59 2621 93
rect 2655 59 2665 93
rect 2603 47 2665 59
rect 2695 161 2749 177
rect 2695 127 2705 161
rect 2739 127 2749 161
rect 2695 93 2749 127
rect 2695 59 2705 93
rect 2739 59 2749 93
rect 2695 47 2749 59
rect 2779 93 2853 177
rect 2779 59 2799 93
rect 2833 59 2853 93
rect 2779 47 2853 59
rect 2883 161 2937 177
rect 2883 127 2893 161
rect 2927 127 2937 161
rect 2883 93 2937 127
rect 2883 59 2893 93
rect 2927 59 2937 93
rect 2883 47 2937 59
rect 2967 93 3019 177
rect 2967 59 2977 93
rect 3011 59 3019 93
rect 3073 135 3125 170
rect 3073 101 3081 135
rect 3115 101 3125 135
rect 3073 66 3125 101
rect 3155 153 3209 170
rect 3155 119 3165 153
rect 3199 119 3209 153
rect 3155 66 3209 119
rect 3239 135 3293 170
rect 3239 101 3249 135
rect 3283 101 3293 135
rect 3239 66 3293 101
rect 3323 153 3377 170
rect 3323 119 3333 153
rect 3367 119 3377 153
rect 3323 66 3377 119
rect 3407 135 3459 170
rect 3407 101 3417 135
rect 3451 101 3459 135
rect 3407 66 3459 101
rect 2967 47 3019 59
rect 3584 106 3636 131
rect 3584 72 3592 106
rect 3626 72 3636 106
rect 3584 47 3636 72
rect 3666 106 3720 131
rect 3666 72 3676 106
rect 3710 72 3720 106
rect 3666 47 3720 72
rect 3750 106 3802 131
rect 3750 72 3760 106
rect 3794 72 3802 106
rect 3750 47 3802 72
rect 3926 106 3978 131
rect 3926 72 3934 106
rect 3968 72 3978 106
rect 3926 47 3978 72
rect 4008 106 4062 131
rect 4008 72 4018 106
rect 4052 72 4062 106
rect 4008 47 4062 72
rect 4092 106 4144 131
rect 4092 72 4102 106
rect 4136 72 4144 106
rect 4092 47 4144 72
rect 4269 135 4321 170
rect 4269 101 4277 135
rect 4311 101 4321 135
rect 4269 66 4321 101
rect 4351 153 4405 170
rect 4351 119 4361 153
rect 4395 119 4405 153
rect 4351 66 4405 119
rect 4435 135 4489 170
rect 4435 101 4445 135
rect 4479 101 4489 135
rect 4435 66 4489 101
rect 4519 153 4573 170
rect 4519 119 4529 153
rect 4563 119 4573 153
rect 4519 66 4573 119
rect 4603 135 4655 170
rect 4603 101 4613 135
rect 4647 101 4655 135
rect 4603 66 4655 101
rect 4709 93 4761 177
rect 4709 59 4717 93
rect 4751 59 4761 93
rect 4709 47 4761 59
rect 4791 161 4845 177
rect 4791 127 4801 161
rect 4835 127 4845 161
rect 4791 93 4845 127
rect 4791 59 4801 93
rect 4835 59 4845 93
rect 4791 47 4845 59
rect 4875 93 4949 177
rect 4875 59 4895 93
rect 4929 59 4949 93
rect 4875 47 4949 59
rect 4979 161 5033 177
rect 4979 127 4989 161
rect 5023 127 5033 161
rect 4979 93 5033 127
rect 4979 59 4989 93
rect 5023 59 5033 93
rect 4979 47 5033 59
rect 5063 161 5125 177
rect 5063 127 5073 161
rect 5107 127 5125 161
rect 5063 93 5125 127
rect 5063 59 5073 93
rect 5107 59 5125 93
rect 5063 47 5125 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 453 497
rect 399 451 411 485
rect 445 451 453 485
rect 998 477 1052 489
rect 399 417 453 451
rect 399 383 411 417
rect 445 383 453 417
rect 399 297 453 383
rect 507 463 561 475
rect 507 429 515 463
rect 549 429 561 463
rect 507 357 561 429
rect 507 323 515 357
rect 549 323 561 357
rect 507 311 561 323
rect 597 425 655 475
rect 597 391 609 425
rect 643 391 655 425
rect 597 357 655 391
rect 597 323 609 357
rect 643 323 655 357
rect 597 311 655 323
rect 691 463 749 475
rect 691 429 703 463
rect 737 429 749 463
rect 691 357 749 429
rect 691 323 703 357
rect 737 323 749 357
rect 691 311 749 323
rect 785 425 843 475
rect 785 391 797 425
rect 831 391 843 425
rect 785 357 843 391
rect 785 323 797 357
rect 831 323 843 357
rect 785 311 843 323
rect 879 463 933 475
rect 879 429 891 463
rect 925 429 933 463
rect 879 363 933 429
rect 879 329 891 363
rect 925 329 933 363
rect 879 311 933 329
rect 998 443 1006 477
rect 1040 443 1052 477
rect 998 371 1052 443
rect 998 337 1006 371
rect 1040 337 1052 371
rect 998 325 1052 337
rect 1088 477 1146 489
rect 1088 443 1100 477
rect 1134 443 1146 477
rect 1088 371 1146 443
rect 1088 337 1100 371
rect 1134 337 1146 371
rect 1088 325 1146 337
rect 1182 477 1236 489
rect 1182 443 1194 477
rect 1228 443 1236 477
rect 1182 371 1236 443
rect 1182 337 1194 371
rect 1228 337 1236 371
rect 1182 325 1236 337
rect 1340 477 1394 489
rect 1340 443 1348 477
rect 1382 443 1394 477
rect 1340 371 1394 443
rect 1340 337 1348 371
rect 1382 337 1394 371
rect 1340 325 1394 337
rect 1430 477 1488 489
rect 1430 443 1442 477
rect 1476 443 1488 477
rect 1430 371 1488 443
rect 1430 337 1442 371
rect 1476 337 1488 371
rect 1430 325 1488 337
rect 1524 477 1578 489
rect 1524 443 1536 477
rect 1570 443 1578 477
rect 2123 485 2177 497
rect 1524 371 1578 443
rect 1524 337 1536 371
rect 1570 337 1578 371
rect 1524 325 1578 337
rect 1643 463 1697 475
rect 1643 429 1651 463
rect 1685 429 1697 463
rect 1643 363 1697 429
rect 1643 329 1651 363
rect 1685 329 1697 363
rect 1643 311 1697 329
rect 1733 425 1791 475
rect 1733 391 1745 425
rect 1779 391 1791 425
rect 1733 357 1791 391
rect 1733 323 1745 357
rect 1779 323 1791 357
rect 1733 311 1791 323
rect 1827 463 1885 475
rect 1827 429 1839 463
rect 1873 429 1885 463
rect 1827 357 1885 429
rect 1827 323 1839 357
rect 1873 323 1885 357
rect 1827 311 1885 323
rect 1921 425 1979 475
rect 1921 391 1933 425
rect 1967 391 1979 425
rect 1921 357 1979 391
rect 1921 323 1933 357
rect 1967 323 1979 357
rect 1921 311 1979 323
rect 2015 463 2069 475
rect 2015 429 2027 463
rect 2061 429 2069 463
rect 2015 357 2069 429
rect 2015 323 2027 357
rect 2061 323 2069 357
rect 2015 311 2069 323
rect 2123 451 2131 485
rect 2165 451 2177 485
rect 2123 417 2177 451
rect 2123 383 2131 417
rect 2165 383 2177 417
rect 2123 297 2177 383
rect 2213 485 2271 497
rect 2213 451 2225 485
rect 2259 451 2271 485
rect 2213 417 2271 451
rect 2213 383 2225 417
rect 2259 383 2271 417
rect 2213 349 2271 383
rect 2213 315 2225 349
rect 2259 315 2271 349
rect 2213 297 2271 315
rect 2307 485 2365 497
rect 2307 451 2319 485
rect 2353 451 2365 485
rect 2307 417 2365 451
rect 2307 383 2319 417
rect 2353 383 2365 417
rect 2307 297 2365 383
rect 2401 485 2459 497
rect 2401 451 2413 485
rect 2447 451 2459 485
rect 2401 417 2459 451
rect 2401 383 2413 417
rect 2447 383 2459 417
rect 2401 349 2459 383
rect 2401 315 2413 349
rect 2447 315 2459 349
rect 2401 297 2459 315
rect 2495 485 2549 497
rect 2495 451 2507 485
rect 2541 451 2549 485
rect 2495 417 2549 451
rect 2495 383 2507 417
rect 2541 383 2549 417
rect 2495 349 2549 383
rect 2495 315 2507 349
rect 2541 315 2549 349
rect 2495 297 2549 315
rect 2603 485 2657 497
rect 2603 451 2611 485
rect 2645 451 2657 485
rect 2603 417 2657 451
rect 2603 383 2611 417
rect 2645 383 2657 417
rect 2603 349 2657 383
rect 2603 315 2611 349
rect 2645 315 2657 349
rect 2603 297 2657 315
rect 2693 485 2751 497
rect 2693 451 2705 485
rect 2739 451 2751 485
rect 2693 417 2751 451
rect 2693 383 2705 417
rect 2739 383 2751 417
rect 2693 349 2751 383
rect 2693 315 2705 349
rect 2739 315 2751 349
rect 2693 297 2751 315
rect 2787 485 2845 497
rect 2787 451 2799 485
rect 2833 451 2845 485
rect 2787 417 2845 451
rect 2787 383 2799 417
rect 2833 383 2845 417
rect 2787 297 2845 383
rect 2881 485 2939 497
rect 2881 451 2893 485
rect 2927 451 2939 485
rect 2881 417 2939 451
rect 2881 383 2893 417
rect 2927 383 2939 417
rect 2881 349 2939 383
rect 2881 315 2893 349
rect 2927 315 2939 349
rect 2881 297 2939 315
rect 2975 485 3029 497
rect 2975 451 2987 485
rect 3021 451 3029 485
rect 3574 477 3628 489
rect 2975 417 3029 451
rect 2975 383 2987 417
rect 3021 383 3029 417
rect 2975 297 3029 383
rect 3083 463 3137 475
rect 3083 429 3091 463
rect 3125 429 3137 463
rect 3083 357 3137 429
rect 3083 323 3091 357
rect 3125 323 3137 357
rect 3083 311 3137 323
rect 3173 425 3231 475
rect 3173 391 3185 425
rect 3219 391 3231 425
rect 3173 357 3231 391
rect 3173 323 3185 357
rect 3219 323 3231 357
rect 3173 311 3231 323
rect 3267 463 3325 475
rect 3267 429 3279 463
rect 3313 429 3325 463
rect 3267 357 3325 429
rect 3267 323 3279 357
rect 3313 323 3325 357
rect 3267 311 3325 323
rect 3361 425 3419 475
rect 3361 391 3373 425
rect 3407 391 3419 425
rect 3361 357 3419 391
rect 3361 323 3373 357
rect 3407 323 3419 357
rect 3361 311 3419 323
rect 3455 463 3509 475
rect 3455 429 3467 463
rect 3501 429 3509 463
rect 3455 363 3509 429
rect 3455 329 3467 363
rect 3501 329 3509 363
rect 3455 311 3509 329
rect 3574 443 3582 477
rect 3616 443 3628 477
rect 3574 371 3628 443
rect 3574 337 3582 371
rect 3616 337 3628 371
rect 3574 325 3628 337
rect 3664 477 3722 489
rect 3664 443 3676 477
rect 3710 443 3722 477
rect 3664 371 3722 443
rect 3664 337 3676 371
rect 3710 337 3722 371
rect 3664 325 3722 337
rect 3758 477 3812 489
rect 3758 443 3770 477
rect 3804 443 3812 477
rect 3758 371 3812 443
rect 3758 337 3770 371
rect 3804 337 3812 371
rect 3758 325 3812 337
rect 3916 477 3970 489
rect 3916 443 3924 477
rect 3958 443 3970 477
rect 3916 371 3970 443
rect 3916 337 3924 371
rect 3958 337 3970 371
rect 3916 325 3970 337
rect 4006 477 4064 489
rect 4006 443 4018 477
rect 4052 443 4064 477
rect 4006 371 4064 443
rect 4006 337 4018 371
rect 4052 337 4064 371
rect 4006 325 4064 337
rect 4100 477 4154 489
rect 4100 443 4112 477
rect 4146 443 4154 477
rect 4699 485 4753 497
rect 4100 371 4154 443
rect 4100 337 4112 371
rect 4146 337 4154 371
rect 4100 325 4154 337
rect 4219 463 4273 475
rect 4219 429 4227 463
rect 4261 429 4273 463
rect 4219 363 4273 429
rect 4219 329 4227 363
rect 4261 329 4273 363
rect 4219 311 4273 329
rect 4309 425 4367 475
rect 4309 391 4321 425
rect 4355 391 4367 425
rect 4309 357 4367 391
rect 4309 323 4321 357
rect 4355 323 4367 357
rect 4309 311 4367 323
rect 4403 463 4461 475
rect 4403 429 4415 463
rect 4449 429 4461 463
rect 4403 357 4461 429
rect 4403 323 4415 357
rect 4449 323 4461 357
rect 4403 311 4461 323
rect 4497 425 4555 475
rect 4497 391 4509 425
rect 4543 391 4555 425
rect 4497 357 4555 391
rect 4497 323 4509 357
rect 4543 323 4555 357
rect 4497 311 4555 323
rect 4591 463 4645 475
rect 4591 429 4603 463
rect 4637 429 4645 463
rect 4591 357 4645 429
rect 4591 323 4603 357
rect 4637 323 4645 357
rect 4591 311 4645 323
rect 4699 451 4707 485
rect 4741 451 4753 485
rect 4699 417 4753 451
rect 4699 383 4707 417
rect 4741 383 4753 417
rect 4699 297 4753 383
rect 4789 485 4847 497
rect 4789 451 4801 485
rect 4835 451 4847 485
rect 4789 417 4847 451
rect 4789 383 4801 417
rect 4835 383 4847 417
rect 4789 349 4847 383
rect 4789 315 4801 349
rect 4835 315 4847 349
rect 4789 297 4847 315
rect 4883 485 4941 497
rect 4883 451 4895 485
rect 4929 451 4941 485
rect 4883 417 4941 451
rect 4883 383 4895 417
rect 4929 383 4941 417
rect 4883 297 4941 383
rect 4977 485 5035 497
rect 4977 451 4989 485
rect 5023 451 5035 485
rect 4977 417 5035 451
rect 4977 383 4989 417
rect 5023 383 5035 417
rect 4977 349 5035 383
rect 4977 315 4989 349
rect 5023 315 5035 349
rect 4977 297 5035 315
rect 5071 485 5125 497
rect 5071 451 5083 485
rect 5117 451 5125 485
rect 5071 417 5125 451
rect 5071 383 5083 417
rect 5117 383 5125 417
rect 5071 349 5125 383
rect 5071 315 5083 349
rect 5117 315 5125 349
rect 5071 297 5125 315
<< ndiffc >>
rect 45 127 79 161
rect 45 59 79 93
rect 129 127 163 161
rect 129 59 163 93
rect 223 59 257 93
rect 317 127 351 161
rect 317 59 351 93
rect 401 59 435 93
rect 505 101 539 135
rect 589 119 623 153
rect 673 101 707 135
rect 757 119 791 153
rect 841 101 875 135
rect 1016 72 1050 106
rect 1100 72 1134 106
rect 1184 72 1218 106
rect 1358 72 1392 106
rect 1442 72 1476 106
rect 1526 72 1560 106
rect 1701 101 1735 135
rect 1785 119 1819 153
rect 1869 101 1903 135
rect 1953 119 1987 153
rect 2037 101 2071 135
rect 2141 59 2175 93
rect 2225 127 2259 161
rect 2225 59 2259 93
rect 2319 59 2353 93
rect 2413 127 2447 161
rect 2413 59 2447 93
rect 2497 127 2531 161
rect 2497 59 2531 93
rect 2621 127 2655 161
rect 2621 59 2655 93
rect 2705 127 2739 161
rect 2705 59 2739 93
rect 2799 59 2833 93
rect 2893 127 2927 161
rect 2893 59 2927 93
rect 2977 59 3011 93
rect 3081 101 3115 135
rect 3165 119 3199 153
rect 3249 101 3283 135
rect 3333 119 3367 153
rect 3417 101 3451 135
rect 3592 72 3626 106
rect 3676 72 3710 106
rect 3760 72 3794 106
rect 3934 72 3968 106
rect 4018 72 4052 106
rect 4102 72 4136 106
rect 4277 101 4311 135
rect 4361 119 4395 153
rect 4445 101 4479 135
rect 4529 119 4563 153
rect 4613 101 4647 135
rect 4717 59 4751 93
rect 4801 127 4835 161
rect 4801 59 4835 93
rect 4895 59 4929 93
rect 4989 127 5023 161
rect 4989 59 5023 93
rect 5073 127 5107 161
rect 5073 59 5107 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 515 429 549 463
rect 515 323 549 357
rect 609 391 643 425
rect 609 323 643 357
rect 703 429 737 463
rect 703 323 737 357
rect 797 391 831 425
rect 797 323 831 357
rect 891 429 925 463
rect 891 329 925 363
rect 1006 443 1040 477
rect 1006 337 1040 371
rect 1100 443 1134 477
rect 1100 337 1134 371
rect 1194 443 1228 477
rect 1194 337 1228 371
rect 1348 443 1382 477
rect 1348 337 1382 371
rect 1442 443 1476 477
rect 1442 337 1476 371
rect 1536 443 1570 477
rect 1536 337 1570 371
rect 1651 429 1685 463
rect 1651 329 1685 363
rect 1745 391 1779 425
rect 1745 323 1779 357
rect 1839 429 1873 463
rect 1839 323 1873 357
rect 1933 391 1967 425
rect 1933 323 1967 357
rect 2027 429 2061 463
rect 2027 323 2061 357
rect 2131 451 2165 485
rect 2131 383 2165 417
rect 2225 451 2259 485
rect 2225 383 2259 417
rect 2225 315 2259 349
rect 2319 451 2353 485
rect 2319 383 2353 417
rect 2413 451 2447 485
rect 2413 383 2447 417
rect 2413 315 2447 349
rect 2507 451 2541 485
rect 2507 383 2541 417
rect 2507 315 2541 349
rect 2611 451 2645 485
rect 2611 383 2645 417
rect 2611 315 2645 349
rect 2705 451 2739 485
rect 2705 383 2739 417
rect 2705 315 2739 349
rect 2799 451 2833 485
rect 2799 383 2833 417
rect 2893 451 2927 485
rect 2893 383 2927 417
rect 2893 315 2927 349
rect 2987 451 3021 485
rect 2987 383 3021 417
rect 3091 429 3125 463
rect 3091 323 3125 357
rect 3185 391 3219 425
rect 3185 323 3219 357
rect 3279 429 3313 463
rect 3279 323 3313 357
rect 3373 391 3407 425
rect 3373 323 3407 357
rect 3467 429 3501 463
rect 3467 329 3501 363
rect 3582 443 3616 477
rect 3582 337 3616 371
rect 3676 443 3710 477
rect 3676 337 3710 371
rect 3770 443 3804 477
rect 3770 337 3804 371
rect 3924 443 3958 477
rect 3924 337 3958 371
rect 4018 443 4052 477
rect 4018 337 4052 371
rect 4112 443 4146 477
rect 4112 337 4146 371
rect 4227 429 4261 463
rect 4227 329 4261 363
rect 4321 391 4355 425
rect 4321 323 4355 357
rect 4415 429 4449 463
rect 4415 323 4449 357
rect 4509 391 4543 425
rect 4509 323 4543 357
rect 4603 429 4637 463
rect 4603 323 4637 357
rect 4707 451 4741 485
rect 4707 383 4741 417
rect 4801 451 4835 485
rect 4801 383 4835 417
rect 4801 315 4835 349
rect 4895 451 4929 485
rect 4895 383 4929 417
rect 4989 451 5023 485
rect 4989 383 5023 417
rect 4989 315 5023 349
rect 5083 451 5117 485
rect 5083 383 5117 417
rect 5083 315 5117 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 561 475 597 523
rect 655 475 691 523
rect 749 475 785 523
rect 843 475 879 523
rect 1052 489 1088 523
rect 1146 489 1182 523
rect 1394 489 1430 523
rect 1488 489 1524 523
rect 1697 475 1733 523
rect 1791 475 1827 523
rect 1885 475 1921 523
rect 1979 475 2015 523
rect 2177 497 2213 523
rect 2271 497 2307 523
rect 2365 497 2401 523
rect 2459 497 2495 523
rect 2657 497 2693 523
rect 2751 497 2787 523
rect 2845 497 2881 523
rect 2939 497 2975 523
rect 81 259 117 297
rect 175 259 211 297
rect 269 259 305 297
rect 363 259 399 297
rect 561 295 597 311
rect 655 295 691 311
rect 749 295 785 311
rect 843 295 879 311
rect 1052 310 1088 325
rect 1146 310 1182 325
rect 1394 310 1430 325
rect 1488 310 1524 325
rect 559 273 925 295
rect 559 265 1008 273
rect 874 263 1008 265
rect 79 249 401 259
rect 79 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 401 249
rect 874 229 890 263
rect 924 229 958 263
rect 992 229 1008 263
rect 874 219 1008 229
rect 79 205 401 215
rect 89 177 119 205
rect 173 177 203 205
rect 277 177 307 205
rect 361 177 391 205
rect 549 170 579 196
rect 633 170 663 196
rect 717 170 747 196
rect 801 170 831 196
rect 1050 177 1090 310
rect 1144 265 1184 310
rect 1392 265 1432 310
rect 1144 249 1267 265
rect 1144 215 1155 249
rect 1189 215 1223 249
rect 1257 215 1267 249
rect 1144 199 1267 215
rect 1309 249 1432 265
rect 1309 215 1319 249
rect 1353 215 1387 249
rect 1421 215 1432 249
rect 1309 199 1432 215
rect 1144 177 1174 199
rect 953 147 1174 177
rect 549 51 579 66
rect 633 51 663 66
rect 717 51 747 66
rect 801 51 831 66
rect 953 51 983 147
rect 1060 131 1090 147
rect 1144 131 1174 147
rect 1402 177 1432 199
rect 1486 177 1526 310
rect 1697 295 1733 311
rect 1791 295 1827 311
rect 1885 295 1921 311
rect 1979 295 2015 311
rect 3137 475 3173 523
rect 3231 475 3267 523
rect 3325 475 3361 523
rect 3419 475 3455 523
rect 3628 489 3664 523
rect 3722 489 3758 523
rect 3970 489 4006 523
rect 4064 489 4100 523
rect 4273 475 4309 523
rect 4367 475 4403 523
rect 4461 475 4497 523
rect 4555 475 4591 523
rect 4753 497 4789 523
rect 4847 497 4883 523
rect 4941 497 4977 523
rect 5035 497 5071 523
rect 1651 273 2017 295
rect 1568 265 2017 273
rect 1568 263 1702 265
rect 1568 229 1584 263
rect 1618 229 1652 263
rect 1686 229 1702 263
rect 2177 259 2213 297
rect 2271 259 2307 297
rect 2365 259 2401 297
rect 2459 259 2495 297
rect 2657 259 2693 297
rect 2751 259 2787 297
rect 2845 259 2881 297
rect 2939 259 2975 297
rect 3137 295 3173 311
rect 3231 295 3267 311
rect 3325 295 3361 311
rect 3419 295 3455 311
rect 3628 310 3664 325
rect 3722 310 3758 325
rect 3970 310 4006 325
rect 4064 310 4100 325
rect 3135 273 3501 295
rect 3135 265 3584 273
rect 3450 263 3584 265
rect 1568 219 1702 229
rect 2175 249 2497 259
rect 2175 215 2235 249
rect 2269 215 2303 249
rect 2337 215 2371 249
rect 2405 215 2439 249
rect 2473 215 2497 249
rect 2175 205 2497 215
rect 2655 249 2977 259
rect 2655 215 2679 249
rect 2713 215 2747 249
rect 2781 215 2815 249
rect 2849 215 2883 249
rect 2917 215 2977 249
rect 3450 229 3466 263
rect 3500 229 3534 263
rect 3568 229 3584 263
rect 3450 219 3584 229
rect 2655 205 2977 215
rect 1402 147 1623 177
rect 1745 170 1775 196
rect 1829 170 1859 196
rect 1913 170 1943 196
rect 1997 170 2027 196
rect 2185 177 2215 205
rect 2269 177 2299 205
rect 2373 177 2403 205
rect 2457 177 2487 205
rect 2665 177 2695 205
rect 2749 177 2779 205
rect 2853 177 2883 205
rect 2937 177 2967 205
rect 1402 131 1432 147
rect 1486 131 1516 147
rect 89 19 119 47
rect 173 21 203 47
rect 277 19 307 47
rect 361 21 391 47
rect 549 21 983 51
rect 1593 51 1623 147
rect 1745 51 1775 66
rect 1829 51 1859 66
rect 1913 51 1943 66
rect 1997 51 2027 66
rect 1060 21 1090 47
rect 1144 21 1174 47
rect 1402 21 1432 47
rect 1486 21 1516 47
rect 1593 21 2027 51
rect 3125 170 3155 196
rect 3209 170 3239 196
rect 3293 170 3323 196
rect 3377 170 3407 196
rect 3626 177 3666 310
rect 3720 265 3760 310
rect 3968 265 4008 310
rect 3720 249 3843 265
rect 3720 215 3731 249
rect 3765 215 3799 249
rect 3833 215 3843 249
rect 3720 199 3843 215
rect 3885 249 4008 265
rect 3885 215 3895 249
rect 3929 215 3963 249
rect 3997 215 4008 249
rect 3885 199 4008 215
rect 3720 177 3750 199
rect 3529 147 3750 177
rect 3125 51 3155 66
rect 3209 51 3239 66
rect 3293 51 3323 66
rect 3377 51 3407 66
rect 3529 51 3559 147
rect 3636 131 3666 147
rect 3720 131 3750 147
rect 3978 177 4008 199
rect 4062 177 4102 310
rect 4273 295 4309 311
rect 4367 295 4403 311
rect 4461 295 4497 311
rect 4555 295 4591 311
rect 4227 273 4593 295
rect 4144 265 4593 273
rect 4144 263 4278 265
rect 4144 229 4160 263
rect 4194 229 4228 263
rect 4262 229 4278 263
rect 4753 259 4789 297
rect 4847 259 4883 297
rect 4941 259 4977 297
rect 5035 259 5071 297
rect 4144 219 4278 229
rect 4751 249 5073 259
rect 4751 215 4811 249
rect 4845 215 4879 249
rect 4913 215 4947 249
rect 4981 215 5015 249
rect 5049 215 5073 249
rect 4751 205 5073 215
rect 3978 147 4199 177
rect 4321 170 4351 196
rect 4405 170 4435 196
rect 4489 170 4519 196
rect 4573 170 4603 196
rect 4761 177 4791 205
rect 4845 177 4875 205
rect 4949 177 4979 205
rect 5033 177 5063 205
rect 3978 131 4008 147
rect 4062 131 4092 147
rect 2185 21 2215 47
rect 2269 19 2299 47
rect 2373 21 2403 47
rect 2457 19 2487 47
rect 2665 19 2695 47
rect 2749 21 2779 47
rect 2853 19 2883 47
rect 2937 21 2967 47
rect 3125 21 3559 51
rect 4169 51 4199 147
rect 4321 51 4351 66
rect 4405 51 4435 66
rect 4489 51 4519 66
rect 4573 51 4603 66
rect 3636 21 3666 47
rect 3720 21 3750 47
rect 3978 21 4008 47
rect 4062 21 4092 47
rect 4169 21 4603 51
rect 4761 21 4791 47
rect 4845 19 4875 47
rect 4949 21 4979 47
rect 5033 19 5063 47
<< polycont >>
rect 103 215 137 249
rect 171 215 205 249
rect 239 215 273 249
rect 307 215 341 249
rect 890 229 924 263
rect 958 229 992 263
rect 1155 215 1189 249
rect 1223 215 1257 249
rect 1319 215 1353 249
rect 1387 215 1421 249
rect 1584 229 1618 263
rect 1652 229 1686 263
rect 2235 215 2269 249
rect 2303 215 2337 249
rect 2371 215 2405 249
rect 2439 215 2473 249
rect 2679 215 2713 249
rect 2747 215 2781 249
rect 2815 215 2849 249
rect 2883 215 2917 249
rect 3466 229 3500 263
rect 3534 229 3568 263
rect 3731 215 3765 249
rect 3799 215 3833 249
rect 3895 215 3929 249
rect 3963 215 3997 249
rect 4160 229 4194 263
rect 4228 229 4262 263
rect 4811 215 4845 249
rect 4879 215 4913 249
rect 4947 215 4981 249
rect 5015 215 5049 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4261 561
rect 4295 527 4353 561
rect 4387 527 4445 561
rect 4479 527 4537 561
rect 4571 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5152 561
rect 25 485 79 527
rect 25 451 35 485
rect 69 451 79 485
rect 25 417 79 451
rect 25 383 35 417
rect 69 383 79 417
rect 25 349 79 383
rect 25 315 35 349
rect 69 315 79 349
rect 25 299 79 315
rect 113 485 179 493
rect 113 451 129 485
rect 163 451 179 485
rect 113 417 179 451
rect 113 383 129 417
rect 163 383 179 417
rect 113 349 179 383
rect 213 485 267 527
rect 213 451 223 485
rect 257 451 267 485
rect 213 417 267 451
rect 213 383 223 417
rect 257 383 267 417
rect 213 367 267 383
rect 301 485 367 493
rect 301 451 317 485
rect 351 451 367 485
rect 301 417 367 451
rect 301 383 317 417
rect 351 383 367 417
rect 113 315 129 349
rect 163 333 179 349
rect 301 349 367 383
rect 401 485 455 527
rect 401 451 411 485
rect 445 451 455 485
rect 401 417 455 451
rect 401 383 411 417
rect 445 383 455 417
rect 401 367 455 383
rect 499 463 941 493
rect 499 429 515 463
rect 549 459 703 463
rect 549 429 559 459
rect 301 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 499 357 559 429
rect 693 429 703 459
rect 737 459 891 463
rect 737 429 747 459
rect 499 333 515 357
rect 351 323 515 333
rect 549 323 559 357
rect 351 315 559 323
rect 113 299 559 315
rect 593 323 609 425
rect 643 323 659 425
rect 593 273 659 323
rect 693 357 747 429
rect 881 429 891 459
rect 925 429 941 463
rect 693 323 703 357
rect 737 323 747 357
rect 693 307 747 323
rect 781 323 797 425
rect 831 323 847 425
rect 781 273 847 323
rect 881 363 941 429
rect 881 329 891 363
rect 925 329 941 363
rect 881 313 941 329
rect 990 477 1045 527
rect 990 443 1006 477
rect 1040 443 1045 477
rect 990 371 1045 443
rect 990 337 1006 371
rect 1040 337 1045 371
rect 990 321 1045 337
rect 1084 477 1150 493
rect 1084 443 1100 477
rect 1134 443 1150 477
rect 1084 371 1150 443
rect 1084 337 1100 371
rect 1134 337 1150 371
rect 1084 321 1150 337
rect 1184 477 1244 527
rect 1184 443 1194 477
rect 1228 443 1244 477
rect 1184 371 1244 443
rect 1184 337 1194 371
rect 1228 337 1244 371
rect 1184 321 1244 337
rect 1332 477 1392 527
rect 1332 443 1348 477
rect 1382 443 1392 477
rect 1332 371 1392 443
rect 1332 337 1348 371
rect 1382 337 1392 371
rect 1332 321 1392 337
rect 1426 477 1492 493
rect 1426 443 1442 477
rect 1476 443 1492 477
rect 1426 371 1492 443
rect 1426 337 1442 371
rect 1476 337 1492 371
rect 1426 321 1492 337
rect 1531 477 1586 527
rect 1531 443 1536 477
rect 1570 443 1586 477
rect 1531 371 1586 443
rect 1531 337 1536 371
rect 1570 337 1586 371
rect 1531 321 1586 337
rect 1635 463 2077 493
rect 1635 429 1651 463
rect 1685 459 1839 463
rect 1685 429 1695 459
rect 1635 363 1695 429
rect 1829 429 1839 459
rect 1873 459 2027 463
rect 1873 429 1883 459
rect 1635 329 1651 363
rect 1685 329 1695 363
rect 1084 279 1118 321
rect 79 249 357 265
rect 79 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 357 249
rect 79 211 357 215
rect 593 213 847 273
rect 881 263 1118 279
rect 1458 279 1492 321
rect 1635 313 1695 329
rect 1729 323 1745 425
rect 1779 323 1795 425
rect 881 229 890 263
rect 924 229 958 263
rect 992 229 1118 263
rect 881 213 1118 229
rect 593 177 639 213
rect 29 161 79 177
rect 29 127 45 161
rect 29 93 79 127
rect 29 59 45 93
rect 29 17 79 59
rect 113 161 539 177
rect 113 127 129 161
rect 163 143 317 161
rect 163 127 179 143
rect 113 93 179 127
rect 301 127 317 143
rect 351 143 539 161
rect 351 127 367 143
rect 113 59 129 93
rect 163 59 179 93
rect 113 51 179 59
rect 213 93 267 109
rect 213 59 223 93
rect 257 59 267 93
rect 213 17 267 59
rect 301 93 367 127
rect 485 135 539 143
rect 301 59 317 93
rect 351 59 367 93
rect 301 51 367 59
rect 401 93 451 109
rect 435 59 451 93
rect 401 17 451 59
rect 485 101 505 135
rect 573 153 639 177
rect 573 119 589 153
rect 623 119 639 153
rect 673 135 707 154
rect 485 85 539 101
rect 741 153 807 213
rect 1084 165 1118 213
rect 1152 249 1271 265
rect 1152 215 1155 249
rect 1189 215 1223 249
rect 1257 215 1271 249
rect 1152 199 1271 215
rect 1305 249 1424 265
rect 1305 215 1319 249
rect 1353 215 1387 249
rect 1421 215 1424 249
rect 1305 199 1424 215
rect 1458 263 1695 279
rect 1458 229 1584 263
rect 1618 229 1652 263
rect 1686 229 1695 263
rect 1458 213 1695 229
rect 1729 273 1795 323
rect 1829 357 1883 429
rect 2017 429 2027 459
rect 2061 429 2077 463
rect 1829 323 1839 357
rect 1873 323 1883 357
rect 1829 307 1883 323
rect 1917 323 1933 425
rect 1967 323 1983 425
rect 1917 273 1983 323
rect 2017 357 2077 429
rect 2121 485 2175 527
rect 2121 451 2131 485
rect 2165 451 2175 485
rect 2121 417 2175 451
rect 2121 383 2131 417
rect 2165 383 2175 417
rect 2121 367 2175 383
rect 2209 485 2275 493
rect 2209 451 2225 485
rect 2259 451 2275 485
rect 2209 417 2275 451
rect 2209 383 2225 417
rect 2259 383 2275 417
rect 2017 323 2027 357
rect 2061 333 2077 357
rect 2209 349 2275 383
rect 2309 485 2363 527
rect 2309 451 2319 485
rect 2353 451 2363 485
rect 2309 417 2363 451
rect 2309 383 2319 417
rect 2353 383 2363 417
rect 2309 367 2363 383
rect 2397 485 2463 493
rect 2397 451 2413 485
rect 2447 451 2463 485
rect 2397 417 2463 451
rect 2397 383 2413 417
rect 2447 383 2463 417
rect 2209 333 2225 349
rect 2061 323 2225 333
rect 2017 315 2225 323
rect 2259 333 2275 349
rect 2397 349 2463 383
rect 2397 333 2413 349
rect 2259 315 2413 333
rect 2447 315 2463 349
rect 2017 299 2463 315
rect 2497 485 2551 527
rect 2497 451 2507 485
rect 2541 451 2551 485
rect 2497 417 2551 451
rect 2497 383 2507 417
rect 2541 383 2551 417
rect 2497 349 2551 383
rect 2497 315 2507 349
rect 2541 315 2551 349
rect 2497 299 2551 315
rect 2601 485 2655 527
rect 2601 451 2611 485
rect 2645 451 2655 485
rect 2601 417 2655 451
rect 2601 383 2611 417
rect 2645 383 2655 417
rect 2601 349 2655 383
rect 2601 315 2611 349
rect 2645 315 2655 349
rect 2601 299 2655 315
rect 2689 485 2755 493
rect 2689 451 2705 485
rect 2739 451 2755 485
rect 2689 417 2755 451
rect 2689 383 2705 417
rect 2739 383 2755 417
rect 2689 349 2755 383
rect 2789 485 2843 527
rect 2789 451 2799 485
rect 2833 451 2843 485
rect 2789 417 2843 451
rect 2789 383 2799 417
rect 2833 383 2843 417
rect 2789 367 2843 383
rect 2877 485 2943 493
rect 2877 451 2893 485
rect 2927 451 2943 485
rect 2877 417 2943 451
rect 2877 383 2893 417
rect 2927 383 2943 417
rect 2689 315 2705 349
rect 2739 333 2755 349
rect 2877 349 2943 383
rect 2977 485 3031 527
rect 2977 451 2987 485
rect 3021 451 3031 485
rect 2977 417 3031 451
rect 2977 383 2987 417
rect 3021 383 3031 417
rect 2977 367 3031 383
rect 3075 463 3517 493
rect 3075 429 3091 463
rect 3125 459 3279 463
rect 3125 429 3135 459
rect 2877 333 2893 349
rect 2739 315 2893 333
rect 2927 333 2943 349
rect 3075 357 3135 429
rect 3269 429 3279 459
rect 3313 459 3467 463
rect 3313 429 3323 459
rect 3075 333 3091 357
rect 2927 323 3091 333
rect 3125 323 3135 357
rect 2927 315 3135 323
rect 2689 299 3135 315
rect 3169 323 3185 425
rect 3219 323 3235 425
rect 1729 213 1983 273
rect 3169 273 3235 323
rect 3269 357 3323 429
rect 3457 429 3467 459
rect 3501 429 3517 463
rect 3269 323 3279 357
rect 3313 323 3323 357
rect 3269 307 3323 323
rect 3357 323 3373 425
rect 3407 323 3423 425
rect 3357 273 3423 323
rect 3457 363 3517 429
rect 3457 329 3467 363
rect 3501 329 3517 363
rect 3457 313 3517 329
rect 3566 477 3621 527
rect 3566 443 3582 477
rect 3616 443 3621 477
rect 3566 371 3621 443
rect 3566 337 3582 371
rect 3616 337 3621 371
rect 3566 321 3621 337
rect 3660 477 3726 493
rect 3660 443 3676 477
rect 3710 443 3726 477
rect 3660 371 3726 443
rect 3660 337 3676 371
rect 3710 337 3726 371
rect 3660 321 3726 337
rect 3760 477 3820 527
rect 3760 443 3770 477
rect 3804 443 3820 477
rect 3760 371 3820 443
rect 3760 337 3770 371
rect 3804 337 3820 371
rect 3760 321 3820 337
rect 3908 477 3968 527
rect 3908 443 3924 477
rect 3958 443 3968 477
rect 3908 371 3968 443
rect 3908 337 3924 371
rect 3958 337 3968 371
rect 3908 321 3968 337
rect 4002 477 4068 493
rect 4002 443 4018 477
rect 4052 443 4068 477
rect 4002 371 4068 443
rect 4002 337 4018 371
rect 4052 337 4068 371
rect 4002 321 4068 337
rect 4107 477 4162 527
rect 4107 443 4112 477
rect 4146 443 4162 477
rect 4107 371 4162 443
rect 4107 337 4112 371
rect 4146 337 4162 371
rect 4107 321 4162 337
rect 4211 463 4653 493
rect 4211 429 4227 463
rect 4261 459 4415 463
rect 4261 429 4271 459
rect 4211 363 4271 429
rect 4405 429 4415 459
rect 4449 459 4603 463
rect 4449 429 4459 459
rect 4211 329 4227 363
rect 4261 329 4271 363
rect 3660 279 3694 321
rect 1458 165 1492 213
rect 741 119 757 153
rect 791 119 807 153
rect 841 135 891 154
rect 673 85 707 101
rect 875 101 891 135
rect 841 85 891 101
rect 485 51 891 85
rect 992 106 1050 122
rect 992 72 1016 106
rect 992 17 1050 72
rect 1084 106 1134 165
rect 1084 72 1100 106
rect 1084 56 1134 72
rect 1176 106 1234 122
rect 1176 72 1184 106
rect 1218 72 1234 106
rect 1176 17 1234 72
rect 1342 106 1400 122
rect 1342 72 1358 106
rect 1392 72 1400 106
rect 1342 17 1400 72
rect 1442 106 1492 165
rect 1685 135 1735 154
rect 1476 72 1492 106
rect 1442 56 1492 72
rect 1526 106 1584 122
rect 1560 72 1584 106
rect 1526 17 1584 72
rect 1685 101 1701 135
rect 1769 153 1835 213
rect 1937 177 1983 213
rect 2219 249 2497 265
rect 2219 215 2235 249
rect 2269 215 2303 249
rect 2337 215 2371 249
rect 2405 215 2439 249
rect 2473 215 2497 249
rect 2219 211 2497 215
rect 2655 249 2933 265
rect 2655 215 2679 249
rect 2713 215 2747 249
rect 2781 215 2815 249
rect 2849 215 2883 249
rect 2917 215 2933 249
rect 2655 211 2933 215
rect 3169 213 3423 273
rect 3457 263 3694 279
rect 4034 279 4068 321
rect 4211 313 4271 329
rect 4305 323 4321 425
rect 4355 323 4371 425
rect 3457 229 3466 263
rect 3500 229 3534 263
rect 3568 229 3694 263
rect 3457 213 3694 229
rect 3169 177 3215 213
rect 1769 119 1785 153
rect 1819 119 1835 153
rect 1869 135 1903 154
rect 1685 85 1735 101
rect 1937 153 2003 177
rect 1937 119 1953 153
rect 1987 119 2003 153
rect 2037 161 2463 177
rect 2037 143 2225 161
rect 2037 135 2091 143
rect 1869 85 1903 101
rect 2071 101 2091 135
rect 2209 127 2225 143
rect 2259 143 2413 161
rect 2259 127 2275 143
rect 2037 85 2091 101
rect 1685 51 2091 85
rect 2125 93 2175 109
rect 2125 59 2141 93
rect 2125 17 2175 59
rect 2209 93 2275 127
rect 2397 127 2413 143
rect 2447 127 2463 161
rect 2209 59 2225 93
rect 2259 59 2275 93
rect 2209 51 2275 59
rect 2309 93 2363 109
rect 2309 59 2319 93
rect 2353 59 2363 93
rect 2309 17 2363 59
rect 2397 93 2463 127
rect 2397 59 2413 93
rect 2447 59 2463 93
rect 2397 51 2463 59
rect 2497 161 2547 177
rect 2531 127 2547 161
rect 2497 93 2547 127
rect 2531 59 2547 93
rect 2497 17 2547 59
rect 2605 161 2655 177
rect 2605 127 2621 161
rect 2605 93 2655 127
rect 2605 59 2621 93
rect 2605 17 2655 59
rect 2689 161 3115 177
rect 2689 127 2705 161
rect 2739 143 2893 161
rect 2739 127 2755 143
rect 2689 93 2755 127
rect 2877 127 2893 143
rect 2927 143 3115 161
rect 2927 127 2943 143
rect 2689 59 2705 93
rect 2739 59 2755 93
rect 2689 51 2755 59
rect 2789 93 2843 109
rect 2789 59 2799 93
rect 2833 59 2843 93
rect 2789 17 2843 59
rect 2877 93 2943 127
rect 3061 135 3115 143
rect 2877 59 2893 93
rect 2927 59 2943 93
rect 2877 51 2943 59
rect 2977 93 3027 109
rect 3011 59 3027 93
rect 2977 17 3027 59
rect 3061 101 3081 135
rect 3149 153 3215 177
rect 3149 119 3165 153
rect 3199 119 3215 153
rect 3249 135 3283 154
rect 3061 85 3115 101
rect 3317 153 3383 213
rect 3660 165 3694 213
rect 3728 249 3847 265
rect 3728 215 3731 249
rect 3765 215 3799 249
rect 3833 215 3847 249
rect 3728 199 3847 215
rect 3881 249 4000 265
rect 3881 215 3895 249
rect 3929 215 3963 249
rect 3997 215 4000 249
rect 3881 199 4000 215
rect 4034 263 4271 279
rect 4034 229 4160 263
rect 4194 229 4228 263
rect 4262 229 4271 263
rect 4034 213 4271 229
rect 4305 273 4371 323
rect 4405 357 4459 429
rect 4593 429 4603 459
rect 4637 429 4653 463
rect 4405 323 4415 357
rect 4449 323 4459 357
rect 4405 307 4459 323
rect 4493 323 4509 425
rect 4543 323 4559 425
rect 4493 273 4559 323
rect 4593 357 4653 429
rect 4697 485 4751 527
rect 4697 451 4707 485
rect 4741 451 4751 485
rect 4697 417 4751 451
rect 4697 383 4707 417
rect 4741 383 4751 417
rect 4697 367 4751 383
rect 4785 485 4851 493
rect 4785 451 4801 485
rect 4835 451 4851 485
rect 4785 417 4851 451
rect 4785 383 4801 417
rect 4835 383 4851 417
rect 4593 323 4603 357
rect 4637 333 4653 357
rect 4785 349 4851 383
rect 4885 485 4939 527
rect 4885 451 4895 485
rect 4929 451 4939 485
rect 4885 417 4939 451
rect 4885 383 4895 417
rect 4929 383 4939 417
rect 4885 367 4939 383
rect 4973 485 5039 493
rect 4973 451 4989 485
rect 5023 451 5039 485
rect 4973 417 5039 451
rect 4973 383 4989 417
rect 5023 383 5039 417
rect 4785 333 4801 349
rect 4637 323 4801 333
rect 4593 315 4801 323
rect 4835 333 4851 349
rect 4973 349 5039 383
rect 4973 333 4989 349
rect 4835 315 4989 333
rect 5023 315 5039 349
rect 4593 299 5039 315
rect 5073 485 5127 527
rect 5073 451 5083 485
rect 5117 451 5127 485
rect 5073 417 5127 451
rect 5073 383 5083 417
rect 5117 383 5127 417
rect 5073 349 5127 383
rect 5073 315 5083 349
rect 5117 315 5127 349
rect 5073 299 5127 315
rect 4305 213 4559 273
rect 4034 165 4068 213
rect 3317 119 3333 153
rect 3367 119 3383 153
rect 3417 135 3467 154
rect 3249 85 3283 101
rect 3451 101 3467 135
rect 3417 85 3467 101
rect 3061 51 3467 85
rect 3568 106 3626 122
rect 3568 72 3592 106
rect 3568 17 3626 72
rect 3660 106 3710 165
rect 3660 72 3676 106
rect 3660 56 3710 72
rect 3752 106 3810 122
rect 3752 72 3760 106
rect 3794 72 3810 106
rect 3752 17 3810 72
rect 3918 106 3976 122
rect 3918 72 3934 106
rect 3968 72 3976 106
rect 3918 17 3976 72
rect 4018 106 4068 165
rect 4261 135 4311 154
rect 4052 72 4068 106
rect 4018 56 4068 72
rect 4102 106 4160 122
rect 4136 72 4160 106
rect 4102 17 4160 72
rect 4261 101 4277 135
rect 4345 153 4411 213
rect 4513 177 4559 213
rect 4795 249 5073 265
rect 4795 215 4811 249
rect 4845 215 4879 249
rect 4913 215 4947 249
rect 4981 215 5015 249
rect 5049 215 5073 249
rect 4795 211 5073 215
rect 4345 119 4361 153
rect 4395 119 4411 153
rect 4445 135 4479 154
rect 4261 85 4311 101
rect 4513 153 4579 177
rect 4513 119 4529 153
rect 4563 119 4579 153
rect 4613 161 5039 177
rect 4613 143 4801 161
rect 4613 135 4667 143
rect 4445 85 4479 101
rect 4647 101 4667 135
rect 4785 127 4801 143
rect 4835 143 4989 161
rect 4835 127 4851 143
rect 4613 85 4667 101
rect 4261 51 4667 85
rect 4701 93 4751 109
rect 4701 59 4717 93
rect 4701 17 4751 59
rect 4785 93 4851 127
rect 4973 127 4989 143
rect 5023 127 5039 161
rect 4785 59 4801 93
rect 4835 59 4851 93
rect 4785 51 4851 59
rect 4885 93 4939 109
rect 4885 59 4895 93
rect 4929 59 4939 93
rect 4885 17 4939 59
rect 4973 93 5039 127
rect 4973 59 4989 93
rect 5023 59 5039 93
rect 4973 51 5039 59
rect 5073 161 5123 177
rect 5107 127 5123 161
rect 5073 93 5123 127
rect 5107 59 5123 93
rect 5073 17 5123 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5152 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3433 527 3467 561
rect 3525 527 3559 561
rect 3617 527 3651 561
rect 3709 527 3743 561
rect 3801 527 3835 561
rect 3893 527 3927 561
rect 3985 527 4019 561
rect 4077 527 4111 561
rect 4169 527 4203 561
rect 4261 527 4295 561
rect 4353 527 4387 561
rect 4445 527 4479 561
rect 4537 527 4571 561
rect 4629 527 4663 561
rect 4721 527 4755 561
rect 4813 527 4847 561
rect 4905 527 4939 561
rect 4997 527 5031 561
rect 5089 527 5123 561
rect 609 357 643 391
rect 797 357 831 391
rect 1745 357 1779 391
rect 1933 357 1967 391
rect 3185 357 3219 391
rect 3373 357 3407 391
rect 4321 357 4355 391
rect 4509 357 4543 391
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
rect 3709 -17 3743 17
rect 3801 -17 3835 17
rect 3893 -17 3927 17
rect 3985 -17 4019 17
rect 4077 -17 4111 17
rect 4169 -17 4203 17
rect 4261 -17 4295 17
rect 4353 -17 4387 17
rect 4445 -17 4479 17
rect 4537 -17 4571 17
rect 4629 -17 4663 17
rect 4721 -17 4755 17
rect 4813 -17 4847 17
rect 4905 -17 4939 17
rect 4997 -17 5031 17
rect 5089 -17 5123 17
<< metal1 >>
rect 0 561 5152 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4261 561
rect 4295 527 4353 561
rect 4387 527 4445 561
rect 4479 527 4537 561
rect 4571 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5152 561
rect 0 496 5152 527
rect 597 391 655 397
rect 597 357 609 391
rect 643 388 655 391
rect 785 391 843 397
rect 785 388 797 391
rect 643 360 797 388
rect 643 357 655 360
rect 597 351 655 357
rect 785 357 797 360
rect 831 388 843 391
rect 1733 391 1791 397
rect 1733 388 1745 391
rect 831 360 1745 388
rect 831 357 843 360
rect 785 351 843 357
rect 1733 357 1745 360
rect 1779 388 1791 391
rect 1921 391 1979 397
rect 1921 388 1933 391
rect 1779 360 1933 388
rect 1779 357 1791 360
rect 1733 351 1791 357
rect 1921 357 1933 360
rect 1967 388 1979 391
rect 3173 391 3231 397
rect 3173 388 3185 391
rect 1967 360 3185 388
rect 1967 357 1979 360
rect 1921 351 1979 357
rect 3173 357 3185 360
rect 3219 388 3231 391
rect 3361 391 3419 397
rect 3361 388 3373 391
rect 3219 360 3373 388
rect 3219 357 3231 360
rect 3173 351 3231 357
rect 3361 357 3373 360
rect 3407 388 3419 391
rect 4309 391 4367 397
rect 4309 388 4321 391
rect 3407 360 4321 388
rect 3407 357 3419 360
rect 3361 351 3419 357
rect 4309 357 4321 360
rect 4355 388 4367 391
rect 4497 391 4555 397
rect 4497 388 4509 391
rect 4355 360 4509 388
rect 4355 357 4367 360
rect 4309 351 4367 357
rect 4497 357 4509 360
rect 4543 357 4555 391
rect 4497 351 4555 357
rect 0 17 5152 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5152 17
rect 0 -48 5152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 muxb4to1_4
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 11 nsew power bidirectional
flabel nwell s 5089 527 5123 561 0 FreeSans 200 180 0 0 VPB
port 11 nsew power bidirectional
flabel nwell s 2605 527 2639 561 0 FreeSans 200 0 0 0 VPB
port 11 nsew power bidirectional
flabel nwell s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPB
port 11 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 10 nsew ground bidirectional
flabel pwell s 5089 -17 5123 17 0 FreeSans 200 180 0 0 VNB
port 10 nsew ground bidirectional
flabel pwell s 2605 -17 2639 17 0 FreeSans 200 0 0 0 VNB
port 10 nsew ground bidirectional
flabel pwell s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VNB
port 10 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 9 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 12 nsew power bidirectional
flabel metal1 s 609 357 643 391 0 FreeSans 200 0 0 0 Z
port 13 nsew signal output
flabel metal1 s 5089 -17 5123 17 0 FreeSans 200 180 0 0 VGND
port 9 nsew ground bidirectional
flabel metal1 s 5089 527 5123 561 0 FreeSans 200 180 0 0 VPWR
port 12 nsew power bidirectional
flabel metal1 s 2605 -17 2639 17 0 FreeSans 200 0 0 0 VGND
port 9 nsew ground bidirectional
flabel metal1 s 2605 527 2639 561 0 FreeSans 200 0 0 0 VPWR
port 12 nsew power bidirectional
flabel metal1 s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VGND
port 9 nsew ground bidirectional
flabel metal1 s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPWR
port 12 nsew power bidirectional
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 S[0]
port 8 nsew signal input
flabel locali s 1317 221 1351 255 0 FreeSans 200 0 0 0 S[1]
port 7 nsew signal input
flabel locali s 2421 221 2455 255 0 FreeSans 200 0 0 0 D[1]
port 3 nsew signal input
flabel locali s 2697 221 2731 256 0 FreeSans 200 0 0 0 D[2]
port 2 nsew signal input
flabel locali s 3801 221 3835 255 0 FreeSans 200 0 0 0 S[2]
port 6 nsew signal input
flabel locali s 3893 221 3927 255 0 FreeSans 200 0 0 0 S[3]
port 5 nsew signal input
flabel locali s 4997 221 5031 255 0 FreeSans 200 0 0 0 D[3]
port 1 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 D[0]
port 4 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 5152 544
string GDS_END 3102408
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 3056922
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
