magic
tech sky130A
magscale 1 2
timestamp 1730626507
<< nwell >>
rect 1944 1394 1960 1639
rect 2036 1073 2052 1318
rect 1760 306 1776 551
rect 2036 230 2052 551
rect 2404 306 2420 551
rect 1944 -15 2052 230
<< viali >>
rect 1109 1651 1143 1685
rect 1720 1651 1754 1685
rect 2030 1651 2064 1685
rect 2640 1651 2674 1685
rect 1289 1195 1323 1229
rect 1208 1027 1242 1061
rect 1376 1027 1410 1061
rect 1526 1027 1560 1061
rect 1616 1027 1650 1061
rect 1802 1027 1836 1061
rect 1891 1027 1925 1061
rect 2127 1027 2161 1061
rect 2480 1027 2514 1061
rect 1653 651 1687 685
rect 1250 563 1284 597
rect 1340 563 1374 597
rect 1482 563 1516 597
rect 1650 563 1684 597
rect 1894 563 1928 597
rect 2170 563 2204 597
rect 2260 563 2294 597
rect 2495 563 2529 597
rect 2848 563 2882 597
rect 1112 -61 1146 -27
rect 1734 -61 1768 -27
rect 2125 -61 2159 -27
rect 2746 -61 2780 -27
<< metal1 >>
rect 1906 1852 1998 1948
rect 2826 1852 3117 1948
rect 1045 1685 1155 1691
rect 1045 1651 1109 1685
rect 1143 1651 1155 1685
rect 1045 1645 1155 1651
rect 1708 1685 2076 1691
rect 1708 1651 1720 1685
rect 1754 1651 2030 1685
rect 2064 1651 2076 1685
rect 1708 1645 2076 1651
rect 2628 1685 2900 1691
rect 2628 1651 2640 1685
rect 2674 1651 2900 1685
rect 2628 1645 2900 1651
rect 972 1308 1078 1404
rect 972 316 1068 1308
rect 1270 1186 1280 1238
rect 1332 1186 1342 1238
rect 1440 1179 1446 1231
rect 1498 1179 1504 1231
rect 1446 1159 1504 1179
rect 1446 1107 1572 1159
rect 1096 1061 1254 1067
rect 1096 1027 1208 1061
rect 1242 1027 1254 1061
rect 1096 1021 1254 1027
rect 1096 603 1142 1021
rect 1357 1018 1367 1070
rect 1419 1018 1429 1070
rect 1514 1061 1572 1107
rect 1985 1067 1995 1070
rect 1514 1027 1526 1061
rect 1560 1027 1572 1061
rect 1514 1021 1572 1027
rect 1604 1061 1848 1067
rect 1604 1027 1616 1061
rect 1650 1027 1802 1061
rect 1836 1027 1848 1061
rect 1604 1021 1848 1027
rect 1879 1061 1995 1067
rect 1879 1027 1891 1061
rect 1925 1027 1995 1061
rect 1879 1021 1995 1027
rect 1985 1018 1995 1021
rect 2047 1067 2057 1070
rect 2854 1067 2900 1645
rect 2047 1061 2173 1067
rect 2047 1027 2127 1061
rect 2161 1027 2173 1061
rect 2047 1021 2173 1027
rect 2468 1061 2900 1067
rect 2468 1027 2480 1061
rect 2514 1027 2900 1061
rect 2468 1021 2900 1027
rect 2047 1018 2057 1021
rect 3021 860 3117 1852
rect 2918 764 3117 860
rect 1641 685 1874 691
rect 1641 651 1653 685
rect 1687 651 1874 685
rect 1641 645 1874 651
rect 1096 597 1296 603
rect 1096 563 1250 597
rect 1284 563 1296 597
rect 1096 557 1296 563
rect 1328 597 1528 603
rect 1328 563 1340 597
rect 1374 563 1482 597
rect 1516 563 1528 597
rect 1328 557 1528 563
rect 1631 554 1641 606
rect 1693 554 1703 606
rect 1828 603 1874 645
rect 1828 597 2216 603
rect 1828 563 1894 597
rect 1928 563 2170 597
rect 2204 563 2216 597
rect 1828 557 2216 563
rect 2248 597 2357 603
rect 2248 563 2260 597
rect 2294 563 2357 597
rect 2248 557 2357 563
rect 2351 551 2357 557
rect 2409 597 2541 603
rect 2409 563 2495 597
rect 2529 563 2541 597
rect 2409 557 2541 563
rect 2836 597 2992 603
rect 2836 563 2848 597
rect 2882 563 2992 597
rect 2836 557 2992 563
rect 2409 551 2415 557
rect 972 220 1078 316
rect 2946 -21 2992 557
rect 978 -27 1158 -21
rect 978 -61 1112 -27
rect 1146 -61 1158 -27
rect 978 -67 1158 -61
rect 1722 -27 2171 -21
rect 1722 -61 1734 -27
rect 1768 -61 2125 -27
rect 2159 -61 2171 -27
rect 1722 -67 2171 -61
rect 2734 -27 2992 -21
rect 2734 -61 2746 -27
rect 2780 -61 2992 -27
rect 2734 -67 2992 -61
rect 3021 -228 3117 764
rect 1906 -324 2090 -228
rect 2918 -324 3117 -228
<< via1 >>
rect 1280 1229 1332 1238
rect 1280 1195 1289 1229
rect 1289 1195 1323 1229
rect 1323 1195 1332 1229
rect 1280 1186 1332 1195
rect 1446 1179 1498 1231
rect 1367 1061 1419 1070
rect 1367 1027 1376 1061
rect 1376 1027 1410 1061
rect 1410 1027 1419 1061
rect 1367 1018 1419 1027
rect 1995 1018 2047 1070
rect 1641 597 1693 606
rect 1641 563 1650 597
rect 1650 563 1684 597
rect 1684 563 1693 597
rect 1641 554 1693 563
rect 2357 551 2409 603
<< metal2 >>
rect 1280 1329 1498 1381
rect 1280 1238 1332 1329
rect 1280 1176 1332 1186
rect 1446 1231 1498 1329
rect 1446 1173 1498 1179
rect 1367 1070 1491 1080
rect 1419 1018 1491 1070
rect 1367 1008 1491 1018
rect 1439 684 1491 1008
rect 1995 1070 2047 1080
rect 1995 836 2047 1018
rect 1406 632 1491 684
rect 1745 789 2047 836
rect 1406 294 1458 632
rect 1641 606 1693 616
rect 1745 606 1797 789
rect 1631 554 1641 606
rect 1693 554 1797 606
rect 2357 603 2409 609
rect 1641 544 1693 554
rect 2357 294 2409 551
rect 1406 242 2409 294
use sky130_fd_sc_hd__nand2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1446 0 1 812
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x2
timestamp 1704896540
transform 1 0 1446 0 -1 812
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1170 0 -1 812
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4
timestamp 1704896540
transform 1 0 1446 0 1 812
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1704896540
transform 1 0 1814 0 -1 812
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1704896540
transform 1 0 1722 0 1 812
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1704896540
transform 1 0 2090 0 -1 812
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2090 0 1 812
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  x9
timestamp 1704896540
transform 1 0 2458 0 -1 812
box -38 -48 498 592
use sky130_fd_sc_hd__inv_8  x10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2826 0 -1 1900
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x11
timestamp 1704896540
transform 1 0 2090 0 1 -276
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x12
timestamp 1704896540
transform -1 0 1906 0 -1 1900
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x13
timestamp 1704896540
transform 1 0 1078 0 1 -276
box -38 -48 866 592
<< labels >>
flabel metal1 1006 784 1006 784 0 FreeSans 1600 0 0 0 vdda
port 0 nsew
flabel metal1 3040 812 3040 812 0 FreeSans 1600 0 0 0 vssa
port 1 nsew
flabel metal1 1124 1039 1124 1039 0 FreeSans 800 0 0 0 in
port 2 nsew
flabel metal1 1017 -54 1017 -54 0 FreeSans 800 0 0 0 clk1
port 3 nsew
flabel metal1 1995 -52 1995 -52 0 FreeSans 800 0 0 0 clkb1
port 4 nsew
flabel metal1 1962 1664 1962 1664 0 FreeSans 800 0 0 0 clkb0
port 5 nsew
flabel metal1 1062 1663 1062 1663 0 FreeSans 800 0 0 0 clk0
port 6 nsew
<< end >>
