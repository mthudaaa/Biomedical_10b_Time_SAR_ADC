magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 2614 582
<< pwell >>
rect 1 199 288 203
rect 1000 199 1576 203
rect 2288 199 2575 203
rect 1 177 469 199
rect 819 177 1757 199
rect 2107 177 2575 199
rect 1 43 2575 177
rect 1 21 288 43
rect 509 21 779 43
rect 1000 21 1576 43
rect 1797 21 2067 43
rect 2288 21 2575 43
rect 29 -17 63 21
rect 1225 -17 1351 21
rect 2513 -17 2547 21
<< scnmos >>
rect 89 47 119 177
rect 173 47 203 177
rect 277 69 307 173
rect 361 69 391 173
rect 587 47 617 151
rect 671 47 701 151
rect 897 69 927 173
rect 981 69 1011 173
rect 1085 47 1115 177
rect 1169 47 1199 177
rect 1377 47 1407 177
rect 1461 47 1491 177
rect 1565 69 1595 173
rect 1649 69 1679 173
rect 1875 47 1905 151
rect 1959 47 1989 151
rect 2185 69 2215 173
rect 2269 69 2299 173
rect 2373 47 2403 177
rect 2457 47 2487 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 280 333 316 497
rect 374 333 410 497
rect 572 297 608 497
rect 680 297 716 497
rect 878 333 914 497
rect 972 333 1008 497
rect 1077 297 1113 497
rect 1171 297 1207 497
rect 1369 297 1405 497
rect 1463 297 1499 497
rect 1568 333 1604 497
rect 1662 333 1698 497
rect 1860 297 1896 497
rect 1968 297 2004 497
rect 2166 333 2202 497
rect 2260 333 2296 497
rect 2365 297 2401 497
rect 2459 297 2495 497
<< ndiff >>
rect 27 161 89 177
rect 27 127 45 161
rect 79 127 89 161
rect 27 93 89 127
rect 27 59 45 93
rect 79 59 89 93
rect 27 47 89 59
rect 119 93 173 177
rect 119 59 129 93
rect 163 59 173 93
rect 119 47 173 59
rect 203 173 262 177
rect 203 169 277 173
rect 203 135 218 169
rect 252 135 277 169
rect 203 101 277 135
rect 203 67 218 101
rect 252 69 277 101
rect 307 153 361 173
rect 307 119 317 153
rect 351 119 361 153
rect 307 69 361 119
rect 391 138 443 173
rect 391 104 401 138
rect 435 104 443 138
rect 391 69 443 104
rect 252 67 262 69
rect 203 47 262 67
rect 1026 173 1085 177
rect 535 116 587 151
rect 535 82 543 116
rect 577 82 587 116
rect 535 47 587 82
rect 617 116 671 151
rect 617 82 627 116
rect 661 82 671 116
rect 617 47 671 82
rect 701 116 753 151
rect 701 82 711 116
rect 745 82 753 116
rect 701 47 753 82
rect 845 138 897 173
rect 845 104 853 138
rect 887 104 897 138
rect 845 69 897 104
rect 927 153 981 173
rect 927 119 937 153
rect 971 119 981 153
rect 927 69 981 119
rect 1011 169 1085 173
rect 1011 135 1036 169
rect 1070 135 1085 169
rect 1011 101 1085 135
rect 1011 69 1036 101
rect 1026 67 1036 69
rect 1070 67 1085 101
rect 1026 47 1085 67
rect 1115 93 1169 177
rect 1115 59 1125 93
rect 1159 59 1169 93
rect 1115 47 1169 59
rect 1199 161 1261 177
rect 1199 127 1209 161
rect 1243 127 1261 161
rect 1199 93 1261 127
rect 1199 59 1209 93
rect 1243 59 1261 93
rect 1199 47 1261 59
rect 1315 161 1377 177
rect 1315 127 1333 161
rect 1367 127 1377 161
rect 1315 93 1377 127
rect 1315 59 1333 93
rect 1367 59 1377 93
rect 1315 47 1377 59
rect 1407 93 1461 177
rect 1407 59 1417 93
rect 1451 59 1461 93
rect 1407 47 1461 59
rect 1491 173 1550 177
rect 1491 169 1565 173
rect 1491 135 1506 169
rect 1540 135 1565 169
rect 1491 101 1565 135
rect 1491 67 1506 101
rect 1540 69 1565 101
rect 1595 153 1649 173
rect 1595 119 1605 153
rect 1639 119 1649 153
rect 1595 69 1649 119
rect 1679 138 1731 173
rect 1679 104 1689 138
rect 1723 104 1731 138
rect 1679 69 1731 104
rect 1540 67 1550 69
rect 1491 47 1550 67
rect 2314 173 2373 177
rect 1823 116 1875 151
rect 1823 82 1831 116
rect 1865 82 1875 116
rect 1823 47 1875 82
rect 1905 116 1959 151
rect 1905 82 1915 116
rect 1949 82 1959 116
rect 1905 47 1959 82
rect 1989 116 2041 151
rect 1989 82 1999 116
rect 2033 82 2041 116
rect 1989 47 2041 82
rect 2133 138 2185 173
rect 2133 104 2141 138
rect 2175 104 2185 138
rect 2133 69 2185 104
rect 2215 153 2269 173
rect 2215 119 2225 153
rect 2259 119 2269 153
rect 2215 69 2269 119
rect 2299 169 2373 173
rect 2299 135 2324 169
rect 2358 135 2373 169
rect 2299 101 2373 135
rect 2299 69 2324 101
rect 2314 67 2324 69
rect 2358 67 2373 101
rect 2314 47 2373 67
rect 2403 93 2457 177
rect 2403 59 2413 93
rect 2447 59 2457 93
rect 2403 47 2457 59
rect 2487 161 2549 177
rect 2487 127 2497 161
rect 2531 127 2549 161
rect 2487 93 2549 127
rect 2487 59 2497 93
rect 2531 59 2549 93
rect 2487 47 2549 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 405 175 451
rect 117 371 129 405
rect 163 371 175 405
rect 117 297 175 371
rect 211 477 280 497
rect 211 443 223 477
rect 257 443 280 477
rect 211 373 280 443
rect 211 339 223 373
rect 257 339 280 373
rect 211 333 280 339
rect 316 421 374 497
rect 316 387 328 421
rect 362 387 374 421
rect 316 333 374 387
rect 410 477 464 497
rect 410 443 422 477
rect 456 443 464 477
rect 410 379 464 443
rect 410 345 422 379
rect 456 345 464 379
rect 410 333 464 345
rect 518 479 572 497
rect 518 445 526 479
rect 560 445 572 479
rect 518 411 572 445
rect 518 377 526 411
rect 560 377 572 411
rect 518 343 572 377
rect 211 297 263 333
rect 518 309 526 343
rect 560 309 572 343
rect 518 297 572 309
rect 608 479 680 497
rect 608 445 627 479
rect 661 445 680 479
rect 608 411 680 445
rect 608 377 627 411
rect 661 377 680 411
rect 608 343 680 377
rect 608 309 627 343
rect 661 309 680 343
rect 608 297 680 309
rect 716 479 770 497
rect 716 445 728 479
rect 762 445 770 479
rect 716 411 770 445
rect 716 377 728 411
rect 762 377 770 411
rect 716 343 770 377
rect 716 309 728 343
rect 762 309 770 343
rect 824 477 878 497
rect 824 443 832 477
rect 866 443 878 477
rect 824 379 878 443
rect 824 345 832 379
rect 866 345 878 379
rect 824 333 878 345
rect 914 421 972 497
rect 914 387 926 421
rect 960 387 972 421
rect 914 333 972 387
rect 1008 477 1077 497
rect 1008 443 1031 477
rect 1065 443 1077 477
rect 1008 373 1077 443
rect 1008 339 1031 373
rect 1065 339 1077 373
rect 1008 333 1077 339
rect 716 297 770 309
rect 1025 297 1077 333
rect 1113 485 1171 497
rect 1113 451 1125 485
rect 1159 451 1171 485
rect 1113 405 1171 451
rect 1113 371 1125 405
rect 1159 371 1171 405
rect 1113 297 1171 371
rect 1207 485 1261 497
rect 1207 451 1219 485
rect 1253 451 1261 485
rect 1207 417 1261 451
rect 1207 383 1219 417
rect 1253 383 1261 417
rect 1207 349 1261 383
rect 1207 315 1219 349
rect 1253 315 1261 349
rect 1207 297 1261 315
rect 1315 485 1369 497
rect 1315 451 1323 485
rect 1357 451 1369 485
rect 1315 417 1369 451
rect 1315 383 1323 417
rect 1357 383 1369 417
rect 1315 349 1369 383
rect 1315 315 1323 349
rect 1357 315 1369 349
rect 1315 297 1369 315
rect 1405 485 1463 497
rect 1405 451 1417 485
rect 1451 451 1463 485
rect 1405 405 1463 451
rect 1405 371 1417 405
rect 1451 371 1463 405
rect 1405 297 1463 371
rect 1499 477 1568 497
rect 1499 443 1511 477
rect 1545 443 1568 477
rect 1499 373 1568 443
rect 1499 339 1511 373
rect 1545 339 1568 373
rect 1499 333 1568 339
rect 1604 421 1662 497
rect 1604 387 1616 421
rect 1650 387 1662 421
rect 1604 333 1662 387
rect 1698 477 1752 497
rect 1698 443 1710 477
rect 1744 443 1752 477
rect 1698 379 1752 443
rect 1698 345 1710 379
rect 1744 345 1752 379
rect 1698 333 1752 345
rect 1806 479 1860 497
rect 1806 445 1814 479
rect 1848 445 1860 479
rect 1806 411 1860 445
rect 1806 377 1814 411
rect 1848 377 1860 411
rect 1806 343 1860 377
rect 1499 297 1551 333
rect 1806 309 1814 343
rect 1848 309 1860 343
rect 1806 297 1860 309
rect 1896 479 1968 497
rect 1896 445 1915 479
rect 1949 445 1968 479
rect 1896 411 1968 445
rect 1896 377 1915 411
rect 1949 377 1968 411
rect 1896 343 1968 377
rect 1896 309 1915 343
rect 1949 309 1968 343
rect 1896 297 1968 309
rect 2004 479 2058 497
rect 2004 445 2016 479
rect 2050 445 2058 479
rect 2004 411 2058 445
rect 2004 377 2016 411
rect 2050 377 2058 411
rect 2004 343 2058 377
rect 2004 309 2016 343
rect 2050 309 2058 343
rect 2112 477 2166 497
rect 2112 443 2120 477
rect 2154 443 2166 477
rect 2112 379 2166 443
rect 2112 345 2120 379
rect 2154 345 2166 379
rect 2112 333 2166 345
rect 2202 421 2260 497
rect 2202 387 2214 421
rect 2248 387 2260 421
rect 2202 333 2260 387
rect 2296 477 2365 497
rect 2296 443 2319 477
rect 2353 443 2365 477
rect 2296 373 2365 443
rect 2296 339 2319 373
rect 2353 339 2365 373
rect 2296 333 2365 339
rect 2004 297 2058 309
rect 2313 297 2365 333
rect 2401 485 2459 497
rect 2401 451 2413 485
rect 2447 451 2459 485
rect 2401 405 2459 451
rect 2401 371 2413 405
rect 2447 371 2459 405
rect 2401 297 2459 371
rect 2495 485 2549 497
rect 2495 451 2507 485
rect 2541 451 2549 485
rect 2495 417 2549 451
rect 2495 383 2507 417
rect 2541 383 2549 417
rect 2495 349 2549 383
rect 2495 315 2507 349
rect 2541 315 2549 349
rect 2495 297 2549 315
<< ndiffc >>
rect 45 127 79 161
rect 45 59 79 93
rect 129 59 163 93
rect 218 135 252 169
rect 218 67 252 101
rect 317 119 351 153
rect 401 104 435 138
rect 543 82 577 116
rect 627 82 661 116
rect 711 82 745 116
rect 853 104 887 138
rect 937 119 971 153
rect 1036 135 1070 169
rect 1036 67 1070 101
rect 1125 59 1159 93
rect 1209 127 1243 161
rect 1209 59 1243 93
rect 1333 127 1367 161
rect 1333 59 1367 93
rect 1417 59 1451 93
rect 1506 135 1540 169
rect 1506 67 1540 101
rect 1605 119 1639 153
rect 1689 104 1723 138
rect 1831 82 1865 116
rect 1915 82 1949 116
rect 1999 82 2033 116
rect 2141 104 2175 138
rect 2225 119 2259 153
rect 2324 135 2358 169
rect 2324 67 2358 101
rect 2413 59 2447 93
rect 2497 127 2531 161
rect 2497 59 2531 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 371 163 405
rect 223 443 257 477
rect 223 339 257 373
rect 328 387 362 421
rect 422 443 456 477
rect 422 345 456 379
rect 526 445 560 479
rect 526 377 560 411
rect 526 309 560 343
rect 627 445 661 479
rect 627 377 661 411
rect 627 309 661 343
rect 728 445 762 479
rect 728 377 762 411
rect 728 309 762 343
rect 832 443 866 477
rect 832 345 866 379
rect 926 387 960 421
rect 1031 443 1065 477
rect 1031 339 1065 373
rect 1125 451 1159 485
rect 1125 371 1159 405
rect 1219 451 1253 485
rect 1219 383 1253 417
rect 1219 315 1253 349
rect 1323 451 1357 485
rect 1323 383 1357 417
rect 1323 315 1357 349
rect 1417 451 1451 485
rect 1417 371 1451 405
rect 1511 443 1545 477
rect 1511 339 1545 373
rect 1616 387 1650 421
rect 1710 443 1744 477
rect 1710 345 1744 379
rect 1814 445 1848 479
rect 1814 377 1848 411
rect 1814 309 1848 343
rect 1915 445 1949 479
rect 1915 377 1949 411
rect 1915 309 1949 343
rect 2016 445 2050 479
rect 2016 377 2050 411
rect 2016 309 2050 343
rect 2120 443 2154 477
rect 2120 345 2154 379
rect 2214 387 2248 421
rect 2319 443 2353 477
rect 2319 339 2353 373
rect 2413 451 2447 485
rect 2413 371 2447 405
rect 2507 451 2541 485
rect 2507 383 2541 417
rect 2507 315 2541 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 280 497 316 523
rect 374 497 410 523
rect 572 497 608 523
rect 680 497 716 523
rect 878 497 914 523
rect 972 497 1008 523
rect 1077 497 1113 523
rect 1171 497 1207 523
rect 1369 497 1405 523
rect 1463 497 1499 523
rect 1568 497 1604 523
rect 1662 497 1698 523
rect 1860 497 1896 523
rect 1968 497 2004 523
rect 2166 497 2202 523
rect 2260 497 2296 523
rect 2365 497 2401 523
rect 2459 497 2495 523
rect 81 259 117 297
rect 175 259 211 297
rect 280 295 316 333
rect 374 295 410 333
rect 278 285 486 295
rect 278 265 436 285
rect 49 249 213 259
rect 49 215 65 249
rect 99 215 133 249
rect 167 215 213 249
rect 420 251 436 265
rect 470 251 486 285
rect 572 282 608 297
rect 680 282 716 297
rect 878 295 914 333
rect 972 295 1008 333
rect 802 285 1010 295
rect 570 265 610 282
rect 678 265 718 282
rect 420 241 486 251
rect 564 249 618 265
rect 49 205 213 215
rect 564 215 574 249
rect 608 215 618 249
rect 89 177 119 205
rect 173 177 203 205
rect 564 199 618 215
rect 670 249 724 265
rect 670 215 680 249
rect 714 215 724 249
rect 802 251 818 285
rect 852 265 1010 285
rect 852 251 868 265
rect 1077 259 1113 297
rect 1171 259 1207 297
rect 1369 259 1405 297
rect 1463 259 1499 297
rect 1568 295 1604 333
rect 1662 295 1698 333
rect 1566 285 1774 295
rect 1566 265 1724 285
rect 802 241 868 251
rect 1075 249 1239 259
rect 670 199 724 215
rect 1075 215 1121 249
rect 1155 215 1189 249
rect 1223 215 1239 249
rect 1075 205 1239 215
rect 1337 249 1501 259
rect 1337 215 1353 249
rect 1387 215 1421 249
rect 1455 215 1501 249
rect 1708 251 1724 265
rect 1758 251 1774 285
rect 1860 282 1896 297
rect 1968 282 2004 297
rect 2166 295 2202 333
rect 2260 295 2296 333
rect 2090 285 2298 295
rect 1858 265 1898 282
rect 1966 265 2006 282
rect 1708 241 1774 251
rect 1852 249 1906 265
rect 1337 205 1501 215
rect 1852 215 1862 249
rect 1896 215 1906 249
rect 277 173 307 199
rect 361 173 391 199
rect 458 169 617 199
rect 277 51 307 69
rect 361 51 391 69
rect 458 51 488 169
rect 587 151 617 169
rect 671 169 830 199
rect 897 173 927 199
rect 981 173 1011 199
rect 1085 177 1115 205
rect 1169 177 1199 205
rect 1377 177 1407 205
rect 1461 177 1491 205
rect 1852 199 1906 215
rect 1958 249 2012 265
rect 1958 215 1968 249
rect 2002 215 2012 249
rect 2090 251 2106 285
rect 2140 265 2298 285
rect 2140 251 2156 265
rect 2365 259 2401 297
rect 2459 259 2495 297
rect 2090 241 2156 251
rect 2363 249 2527 259
rect 1958 199 2012 215
rect 2363 215 2409 249
rect 2443 215 2477 249
rect 2511 215 2527 249
rect 2363 205 2527 215
rect 671 151 701 169
rect 89 19 119 47
rect 173 21 203 47
rect 277 21 488 51
rect 800 51 830 169
rect 897 51 927 69
rect 981 51 1011 69
rect 587 21 617 47
rect 671 21 701 47
rect 800 21 1011 51
rect 1565 173 1595 199
rect 1649 173 1679 199
rect 1746 169 1905 199
rect 1565 51 1595 69
rect 1649 51 1679 69
rect 1746 51 1776 169
rect 1875 151 1905 169
rect 1959 169 2118 199
rect 2185 173 2215 199
rect 2269 173 2299 199
rect 2373 177 2403 205
rect 2457 177 2487 205
rect 1959 151 1989 169
rect 1085 21 1115 47
rect 1169 19 1199 47
rect 1377 19 1407 47
rect 1461 21 1491 47
rect 1565 21 1776 51
rect 2088 51 2118 169
rect 2185 51 2215 69
rect 2269 51 2299 69
rect 1875 21 1905 47
rect 1959 21 1989 47
rect 2088 21 2299 51
rect 2373 21 2403 47
rect 2457 19 2487 47
<< polycont >>
rect 65 215 99 249
rect 133 215 167 249
rect 436 251 470 285
rect 574 215 608 249
rect 680 215 714 249
rect 818 251 852 285
rect 1121 215 1155 249
rect 1189 215 1223 249
rect 1353 215 1387 249
rect 1421 215 1455 249
rect 1724 251 1758 285
rect 1862 215 1896 249
rect 1968 215 2002 249
rect 2106 251 2140 285
rect 2409 215 2443 249
rect 2477 215 2511 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 19 485 85 493
rect 19 451 35 485
rect 69 451 85 485
rect 19 442 85 451
rect 119 485 179 527
rect 119 451 129 485
rect 163 451 179 485
rect 19 417 79 442
rect 119 421 179 451
rect 19 383 35 417
rect 69 383 79 417
rect 19 349 79 383
rect 113 405 179 421
rect 113 371 129 405
rect 163 371 179 405
rect 113 367 179 371
rect 223 477 456 493
rect 257 459 422 477
rect 223 373 257 443
rect 19 315 35 349
rect 69 333 79 349
rect 293 421 379 425
rect 293 391 328 421
rect 293 357 305 391
rect 362 387 379 421
rect 339 357 379 387
rect 293 351 379 357
rect 422 379 456 443
rect 223 333 257 339
rect 69 315 257 333
rect 19 299 257 315
rect 19 249 183 265
rect 19 215 65 249
rect 99 215 133 249
rect 167 215 183 249
rect 19 211 183 215
rect 206 177 267 185
rect 317 177 351 351
rect 422 329 456 345
rect 510 479 576 493
rect 510 445 526 479
rect 560 445 576 479
rect 510 411 576 445
rect 510 377 526 411
rect 560 377 576 411
rect 510 343 576 377
rect 510 327 526 343
rect 490 309 526 327
rect 560 309 576 343
rect 490 295 576 309
rect 420 293 576 295
rect 611 479 677 527
rect 611 445 627 479
rect 661 445 677 479
rect 611 411 677 445
rect 611 377 627 411
rect 661 377 677 411
rect 611 343 677 377
rect 611 309 627 343
rect 661 309 677 343
rect 611 293 677 309
rect 712 479 778 493
rect 712 445 728 479
rect 762 445 778 479
rect 712 411 778 445
rect 712 377 728 411
rect 762 377 778 411
rect 712 343 778 377
rect 712 309 728 343
rect 762 327 778 343
rect 832 477 1065 493
rect 866 459 1031 477
rect 832 379 866 443
rect 909 421 995 425
rect 909 387 926 421
rect 960 391 995 421
rect 909 357 949 387
rect 983 357 995 391
rect 909 351 995 357
rect 1031 373 1065 443
rect 832 329 866 345
rect 762 309 798 327
rect 712 295 798 309
rect 712 293 868 295
rect 420 285 524 293
rect 420 251 436 285
rect 470 261 524 285
rect 764 285 868 293
rect 764 261 818 285
rect 470 251 503 261
rect 420 241 503 251
rect 29 169 267 177
rect 29 161 218 169
rect 29 127 45 161
rect 79 143 218 161
rect 79 127 95 143
rect 29 93 95 127
rect 206 135 218 143
rect 252 135 267 169
rect 29 59 45 93
rect 79 59 95 93
rect 29 51 95 59
rect 129 93 172 109
rect 163 59 172 93
rect 129 17 172 59
rect 206 101 267 135
rect 301 153 367 177
rect 301 119 317 153
rect 351 119 367 153
rect 401 138 435 154
rect 206 67 218 101
rect 252 85 267 101
rect 469 151 503 241
rect 558 249 625 259
rect 558 215 574 249
rect 608 215 625 249
rect 558 205 625 215
rect 663 249 730 259
rect 663 215 680 249
rect 714 215 730 249
rect 663 205 730 215
rect 785 251 818 261
rect 852 251 868 285
rect 785 241 868 251
rect 785 151 819 241
rect 937 177 971 351
rect 1109 485 1169 527
rect 1109 451 1125 485
rect 1159 451 1169 485
rect 1109 421 1169 451
rect 1203 485 1269 493
rect 1203 451 1219 485
rect 1253 451 1269 485
rect 1203 442 1269 451
rect 1109 405 1175 421
rect 1109 371 1125 405
rect 1159 371 1175 405
rect 1109 367 1175 371
rect 1209 417 1269 442
rect 1209 383 1219 417
rect 1253 383 1269 417
rect 1031 333 1065 339
rect 1209 349 1269 383
rect 1209 333 1219 349
rect 1031 315 1219 333
rect 1253 315 1269 349
rect 1031 299 1269 315
rect 1307 485 1373 493
rect 1307 451 1323 485
rect 1357 451 1373 485
rect 1307 442 1373 451
rect 1407 485 1467 527
rect 1407 451 1417 485
rect 1451 451 1467 485
rect 1307 417 1367 442
rect 1407 421 1467 451
rect 1307 383 1323 417
rect 1357 383 1367 417
rect 1307 349 1367 383
rect 1401 405 1467 421
rect 1401 371 1417 405
rect 1451 371 1467 405
rect 1401 367 1467 371
rect 1511 477 1744 493
rect 1545 459 1710 477
rect 1511 373 1545 443
rect 1307 315 1323 349
rect 1357 333 1367 349
rect 1581 421 1667 425
rect 1581 391 1616 421
rect 1581 357 1593 391
rect 1650 387 1667 421
rect 1627 357 1667 387
rect 1581 351 1667 357
rect 1710 379 1744 443
rect 1511 333 1545 339
rect 1357 315 1545 333
rect 1307 299 1545 315
rect 1105 249 1269 265
rect 1105 215 1121 249
rect 1155 215 1189 249
rect 1223 215 1269 249
rect 1105 211 1269 215
rect 1307 249 1471 265
rect 1307 215 1353 249
rect 1387 215 1421 249
rect 1455 215 1471 249
rect 1307 211 1471 215
rect 1021 177 1082 185
rect 1494 177 1555 185
rect 1605 177 1639 351
rect 1710 329 1744 345
rect 1798 479 1864 493
rect 1798 445 1814 479
rect 1848 445 1864 479
rect 1798 411 1864 445
rect 1798 377 1814 411
rect 1848 377 1864 411
rect 1798 343 1864 377
rect 1798 327 1814 343
rect 1778 309 1814 327
rect 1848 309 1864 343
rect 1778 295 1864 309
rect 1708 293 1864 295
rect 1899 479 1965 527
rect 1899 445 1915 479
rect 1949 445 1965 479
rect 1899 411 1965 445
rect 1899 377 1915 411
rect 1949 377 1965 411
rect 1899 343 1965 377
rect 1899 309 1915 343
rect 1949 309 1965 343
rect 1899 293 1965 309
rect 2000 479 2066 493
rect 2000 445 2016 479
rect 2050 445 2066 479
rect 2000 411 2066 445
rect 2000 377 2016 411
rect 2050 377 2066 411
rect 2000 343 2066 377
rect 2000 309 2016 343
rect 2050 327 2066 343
rect 2120 477 2353 493
rect 2154 459 2319 477
rect 2120 379 2154 443
rect 2197 421 2283 425
rect 2197 387 2214 421
rect 2248 391 2283 421
rect 2197 357 2237 387
rect 2271 357 2283 391
rect 2197 351 2283 357
rect 2319 373 2353 443
rect 2120 329 2154 345
rect 2050 309 2086 327
rect 2000 295 2086 309
rect 2000 293 2156 295
rect 1708 285 1812 293
rect 1708 251 1724 285
rect 1758 261 1812 285
rect 2052 285 2156 293
rect 2052 261 2106 285
rect 1758 251 1791 261
rect 1708 241 1791 251
rect 469 117 585 151
rect 401 85 435 104
rect 252 67 435 85
rect 206 51 435 67
rect 535 116 585 117
rect 535 82 543 116
rect 577 82 585 116
rect 535 66 585 82
rect 619 116 669 132
rect 619 82 627 116
rect 661 82 669 116
rect 619 17 669 82
rect 703 117 819 151
rect 853 138 887 154
rect 703 116 753 117
rect 703 82 711 116
rect 745 82 753 116
rect 703 66 753 82
rect 921 153 987 177
rect 921 119 937 153
rect 971 119 987 153
rect 1021 169 1259 177
rect 1021 135 1036 169
rect 1070 161 1259 169
rect 1070 143 1209 161
rect 1070 135 1082 143
rect 853 85 887 104
rect 1021 101 1082 135
rect 1193 127 1209 143
rect 1243 127 1259 161
rect 1021 85 1036 101
rect 853 67 1036 85
rect 1070 67 1082 101
rect 853 51 1082 67
rect 1116 93 1159 109
rect 1116 59 1125 93
rect 1116 17 1159 59
rect 1193 93 1259 127
rect 1193 59 1209 93
rect 1243 59 1259 93
rect 1193 51 1259 59
rect 1317 169 1555 177
rect 1317 161 1506 169
rect 1317 127 1333 161
rect 1367 143 1506 161
rect 1367 127 1383 143
rect 1317 93 1383 127
rect 1494 135 1506 143
rect 1540 135 1555 169
rect 1317 59 1333 93
rect 1367 59 1383 93
rect 1317 51 1383 59
rect 1417 93 1460 109
rect 1451 59 1460 93
rect 1417 17 1460 59
rect 1494 101 1555 135
rect 1589 153 1655 177
rect 1589 119 1605 153
rect 1639 119 1655 153
rect 1689 138 1723 154
rect 1494 67 1506 101
rect 1540 85 1555 101
rect 1757 151 1791 241
rect 1846 249 1913 259
rect 1846 215 1862 249
rect 1896 215 1913 249
rect 1846 205 1913 215
rect 1951 249 2018 259
rect 1951 215 1968 249
rect 2002 215 2018 249
rect 1951 205 2018 215
rect 2073 251 2106 261
rect 2140 251 2156 285
rect 2073 241 2156 251
rect 2073 151 2107 241
rect 2225 177 2259 351
rect 2397 485 2457 527
rect 2397 451 2413 485
rect 2447 451 2457 485
rect 2397 421 2457 451
rect 2491 485 2557 493
rect 2491 451 2507 485
rect 2541 451 2557 485
rect 2491 442 2557 451
rect 2397 405 2463 421
rect 2397 371 2413 405
rect 2447 371 2463 405
rect 2397 367 2463 371
rect 2497 417 2557 442
rect 2497 383 2507 417
rect 2541 383 2557 417
rect 2319 333 2353 339
rect 2497 349 2557 383
rect 2497 333 2507 349
rect 2319 315 2507 333
rect 2541 315 2557 349
rect 2319 299 2557 315
rect 2393 249 2557 265
rect 2393 215 2409 249
rect 2443 215 2477 249
rect 2511 215 2557 249
rect 2393 211 2557 215
rect 2309 177 2370 185
rect 1757 117 1873 151
rect 1689 85 1723 104
rect 1540 67 1723 85
rect 1494 51 1723 67
rect 1823 116 1873 117
rect 1823 82 1831 116
rect 1865 82 1873 116
rect 1823 66 1873 82
rect 1907 116 1957 132
rect 1907 82 1915 116
rect 1949 82 1957 116
rect 1907 17 1957 82
rect 1991 117 2107 151
rect 2141 138 2175 154
rect 1991 116 2041 117
rect 1991 82 1999 116
rect 2033 82 2041 116
rect 1991 66 2041 82
rect 2209 153 2275 177
rect 2209 119 2225 153
rect 2259 119 2275 153
rect 2309 169 2547 177
rect 2309 135 2324 169
rect 2358 161 2547 169
rect 2358 143 2497 161
rect 2358 135 2370 143
rect 2141 85 2175 104
rect 2309 101 2370 135
rect 2481 127 2497 143
rect 2531 127 2547 161
rect 2309 85 2324 101
rect 2141 67 2324 85
rect 2358 67 2370 101
rect 2141 51 2370 67
rect 2404 93 2447 109
rect 2404 59 2413 93
rect 2404 17 2447 59
rect 2481 93 2547 127
rect 2481 59 2497 93
rect 2531 59 2547 93
rect 2481 51 2547 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 305 387 328 391
rect 328 387 339 391
rect 305 357 339 387
rect 949 387 960 391
rect 960 387 983 391
rect 949 357 983 387
rect 1593 387 1616 391
rect 1616 387 1627 391
rect 1593 357 1627 387
rect 2237 387 2248 391
rect 2248 387 2271 391
rect 2237 357 2271 387
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
<< metal1 >>
rect 0 561 2576 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 0 496 2576 527
rect 293 391 351 397
rect 293 357 305 391
rect 339 388 351 391
rect 937 391 995 397
rect 937 388 949 391
rect 339 360 949 388
rect 339 357 351 360
rect 293 351 351 357
rect 937 357 949 360
rect 983 388 995 391
rect 1581 391 1639 397
rect 1581 388 1593 391
rect 983 360 1593 388
rect 983 357 995 360
rect 937 351 995 357
rect 1581 357 1593 360
rect 1627 388 1639 391
rect 2225 391 2283 397
rect 2225 388 2237 391
rect 1627 360 2237 388
rect 1627 357 1639 360
rect 1581 351 1639 357
rect 2225 357 2237 360
rect 2271 357 2283 391
rect 2225 351 2283 357
rect 0 17 2576 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
rect 0 -48 2576 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 9 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 12 nsew power bidirectional
flabel metal1 s 305 357 339 391 0 FreeSans 200 0 0 0 Z
port 13 nsew signal output
flabel metal1 s 1317 -17 1351 17 0 FreeSans 200 0 0 0 VGND
port 9 nsew ground bidirectional
flabel metal1 s 1317 527 1351 561 0 FreeSans 200 0 0 0 VPWR
port 12 nsew power bidirectional
flabel metal1 s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPWR
port 12 nsew power bidirectional
flabel metal1 s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VGND
port 9 nsew ground bidirectional
flabel metal1 s 1225 -17 1259 17 0 FreeSans 200 180 0 0 VGND
port 9 nsew ground bidirectional
flabel metal1 s 1225 527 1259 561 0 FreeSans 200 180 0 0 VPWR
port 12 nsew power bidirectional
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 10 nsew ground bidirectional
flabel pwell s 1317 -17 1351 17 0 FreeSans 200 0 0 0 VNB
port 10 nsew ground bidirectional
flabel pwell s 2513 -17 2547 17 0 FreeSans 200 180 0 0 VNB
port 10 nsew ground bidirectional
flabel pwell s 1225 -17 1259 17 0 FreeSans 200 180 0 0 VNB
port 10 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 11 nsew power bidirectional
flabel nwell s 1317 527 1351 561 0 FreeSans 200 0 0 0 VPB
port 11 nsew power bidirectional
flabel nwell s 2513 527 2547 561 0 FreeSans 200 180 0 0 VPB
port 11 nsew power bidirectional
flabel nwell s 1225 527 1259 561 0 FreeSans 200 180 0 0 VPB
port 11 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 muxb4to1_2
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 S[1]
port 7 nsew signal input
flabel locali s 1869 221 1903 255 0 FreeSans 200 0 0 0 S[2]
port 6 nsew signal input
flabel locali s 1961 221 1995 255 0 FreeSans 200 0 0 0 S[3]
port 5 nsew signal input
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 D[1]
port 3 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 D[0]
port 4 nsew signal input
flabel locali s 1317 221 1351 256 0 FreeSans 200 0 0 0 D[2]
port 2 nsew signal input
flabel locali s 2513 221 2547 255 0 FreeSans 200 0 0 0 D[3]
port 1 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 S[0]
port 8 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 2576 544
string GDS_END 3132212
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 3102470
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
