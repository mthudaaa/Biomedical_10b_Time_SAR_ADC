magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 2430 582
<< pwell >>
rect 1 21 2359 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 183 47 213 177
rect 267 47 297 177
rect 371 47 401 177
rect 455 47 485 177
rect 559 47 589 177
rect 643 47 673 177
rect 747 47 777 177
rect 831 47 861 177
rect 935 47 965 177
rect 1019 47 1049 177
rect 1123 47 1153 177
rect 1207 47 1237 177
rect 1301 47 1331 177
rect 1395 47 1425 177
rect 1499 47 1529 177
rect 1583 47 1613 177
rect 1687 47 1717 177
rect 1771 47 1801 177
rect 1865 47 1895 177
rect 1959 47 1989 177
rect 2063 47 2093 177
rect 2147 47 2177 177
rect 2251 47 2281 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
rect 1209 297 1245 497
rect 1303 297 1339 497
rect 1397 297 1433 497
rect 1491 297 1527 497
rect 1585 297 1621 497
rect 1679 297 1715 497
rect 1773 297 1809 497
rect 1867 297 1903 497
rect 1961 297 1997 497
rect 2055 297 2091 497
rect 2149 297 2185 497
rect 2243 297 2279 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 93 183 177
rect 109 59 129 93
rect 163 59 183 93
rect 109 47 183 59
rect 213 161 267 177
rect 213 127 223 161
rect 257 127 267 161
rect 213 93 267 127
rect 213 59 223 93
rect 257 59 267 93
rect 213 47 267 59
rect 297 93 371 177
rect 297 59 317 93
rect 351 59 371 93
rect 297 47 371 59
rect 401 161 455 177
rect 401 127 411 161
rect 445 127 455 161
rect 401 93 455 127
rect 401 59 411 93
rect 445 59 455 93
rect 401 47 455 59
rect 485 93 559 177
rect 485 59 505 93
rect 539 59 559 93
rect 485 47 559 59
rect 589 161 643 177
rect 589 127 599 161
rect 633 127 643 161
rect 589 93 643 127
rect 589 59 599 93
rect 633 59 643 93
rect 589 47 643 59
rect 673 93 747 177
rect 673 59 693 93
rect 727 59 747 93
rect 673 47 747 59
rect 777 161 831 177
rect 777 127 787 161
rect 821 127 831 161
rect 777 93 831 127
rect 777 59 787 93
rect 821 59 831 93
rect 777 47 831 59
rect 861 93 935 177
rect 861 59 881 93
rect 915 59 935 93
rect 861 47 935 59
rect 965 161 1019 177
rect 965 127 975 161
rect 1009 127 1019 161
rect 965 93 1019 127
rect 965 59 975 93
rect 1009 59 1019 93
rect 965 47 1019 59
rect 1049 93 1123 177
rect 1049 59 1069 93
rect 1103 59 1123 93
rect 1049 47 1123 59
rect 1153 161 1207 177
rect 1153 127 1163 161
rect 1197 127 1207 161
rect 1153 93 1207 127
rect 1153 59 1163 93
rect 1197 59 1207 93
rect 1153 47 1207 59
rect 1237 161 1301 177
rect 1237 127 1257 161
rect 1291 127 1301 161
rect 1237 47 1301 127
rect 1331 93 1395 177
rect 1331 59 1351 93
rect 1385 59 1395 93
rect 1331 47 1395 59
rect 1425 161 1499 177
rect 1425 127 1445 161
rect 1479 127 1499 161
rect 1425 47 1499 127
rect 1529 93 1583 177
rect 1529 59 1539 93
rect 1573 59 1583 93
rect 1529 47 1583 59
rect 1613 161 1687 177
rect 1613 127 1633 161
rect 1667 127 1687 161
rect 1613 47 1687 127
rect 1717 93 1771 177
rect 1717 59 1727 93
rect 1761 59 1771 93
rect 1717 47 1771 59
rect 1801 161 1865 177
rect 1801 127 1821 161
rect 1855 127 1865 161
rect 1801 47 1865 127
rect 1895 93 1959 177
rect 1895 59 1915 93
rect 1949 59 1959 93
rect 1895 47 1959 59
rect 1989 161 2063 177
rect 1989 127 2009 161
rect 2043 127 2063 161
rect 1989 47 2063 127
rect 2093 93 2147 177
rect 2093 59 2103 93
rect 2137 59 2147 93
rect 2093 47 2147 59
rect 2177 161 2251 177
rect 2177 127 2197 161
rect 2231 127 2251 161
rect 2177 47 2251 127
rect 2281 161 2333 177
rect 2281 127 2291 161
rect 2325 127 2333 161
rect 2281 93 2333 127
rect 2281 59 2291 93
rect 2325 59 2333 93
rect 2281 47 2333 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 349 551 383
rect 493 315 505 349
rect 539 315 551 349
rect 493 297 551 315
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 417 645 451
rect 587 383 599 417
rect 633 383 645 417
rect 587 297 645 383
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 349 739 383
rect 681 315 693 349
rect 727 315 739 349
rect 681 297 739 315
rect 775 485 833 497
rect 775 451 787 485
rect 821 451 833 485
rect 775 417 833 451
rect 775 383 787 417
rect 821 383 833 417
rect 775 297 833 383
rect 869 485 927 497
rect 869 451 881 485
rect 915 451 927 485
rect 869 417 927 451
rect 869 383 881 417
rect 915 383 927 417
rect 869 349 927 383
rect 869 315 881 349
rect 915 315 927 349
rect 869 297 927 315
rect 963 485 1021 497
rect 963 451 975 485
rect 1009 451 1021 485
rect 963 417 1021 451
rect 963 383 975 417
rect 1009 383 1021 417
rect 963 297 1021 383
rect 1057 485 1115 497
rect 1057 451 1069 485
rect 1103 451 1115 485
rect 1057 417 1115 451
rect 1057 383 1069 417
rect 1103 383 1115 417
rect 1057 349 1115 383
rect 1057 315 1069 349
rect 1103 315 1115 349
rect 1057 297 1115 315
rect 1151 485 1209 497
rect 1151 451 1163 485
rect 1197 451 1209 485
rect 1151 417 1209 451
rect 1151 383 1163 417
rect 1197 383 1209 417
rect 1151 297 1209 383
rect 1245 485 1303 497
rect 1245 451 1257 485
rect 1291 451 1303 485
rect 1245 417 1303 451
rect 1245 383 1257 417
rect 1291 383 1303 417
rect 1245 349 1303 383
rect 1245 315 1257 349
rect 1291 315 1303 349
rect 1245 297 1303 315
rect 1339 485 1397 497
rect 1339 451 1351 485
rect 1385 451 1397 485
rect 1339 417 1397 451
rect 1339 383 1351 417
rect 1385 383 1397 417
rect 1339 297 1397 383
rect 1433 485 1491 497
rect 1433 451 1445 485
rect 1479 451 1491 485
rect 1433 417 1491 451
rect 1433 383 1445 417
rect 1479 383 1491 417
rect 1433 349 1491 383
rect 1433 315 1445 349
rect 1479 315 1491 349
rect 1433 297 1491 315
rect 1527 485 1585 497
rect 1527 451 1539 485
rect 1573 451 1585 485
rect 1527 417 1585 451
rect 1527 383 1539 417
rect 1573 383 1585 417
rect 1527 297 1585 383
rect 1621 485 1679 497
rect 1621 451 1633 485
rect 1667 451 1679 485
rect 1621 417 1679 451
rect 1621 383 1633 417
rect 1667 383 1679 417
rect 1621 349 1679 383
rect 1621 315 1633 349
rect 1667 315 1679 349
rect 1621 297 1679 315
rect 1715 485 1773 497
rect 1715 451 1727 485
rect 1761 451 1773 485
rect 1715 417 1773 451
rect 1715 383 1727 417
rect 1761 383 1773 417
rect 1715 297 1773 383
rect 1809 485 1867 497
rect 1809 451 1821 485
rect 1855 451 1867 485
rect 1809 417 1867 451
rect 1809 383 1821 417
rect 1855 383 1867 417
rect 1809 349 1867 383
rect 1809 315 1821 349
rect 1855 315 1867 349
rect 1809 297 1867 315
rect 1903 485 1961 497
rect 1903 451 1915 485
rect 1949 451 1961 485
rect 1903 417 1961 451
rect 1903 383 1915 417
rect 1949 383 1961 417
rect 1903 297 1961 383
rect 1997 485 2055 497
rect 1997 451 2009 485
rect 2043 451 2055 485
rect 1997 417 2055 451
rect 1997 383 2009 417
rect 2043 383 2055 417
rect 1997 349 2055 383
rect 1997 315 2009 349
rect 2043 315 2055 349
rect 1997 297 2055 315
rect 2091 485 2149 497
rect 2091 451 2103 485
rect 2137 451 2149 485
rect 2091 417 2149 451
rect 2091 383 2103 417
rect 2137 383 2149 417
rect 2091 297 2149 383
rect 2185 485 2243 497
rect 2185 451 2197 485
rect 2231 451 2243 485
rect 2185 417 2243 451
rect 2185 383 2197 417
rect 2231 383 2243 417
rect 2185 349 2243 383
rect 2185 315 2197 349
rect 2231 315 2243 349
rect 2185 297 2243 315
rect 2279 485 2333 497
rect 2279 451 2291 485
rect 2325 451 2333 485
rect 2279 417 2333 451
rect 2279 383 2291 417
rect 2325 383 2333 417
rect 2279 349 2333 383
rect 2279 315 2291 349
rect 2325 315 2333 349
rect 2279 297 2333 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 59 163 93
rect 223 127 257 161
rect 223 59 257 93
rect 317 59 351 93
rect 411 127 445 161
rect 411 59 445 93
rect 505 59 539 93
rect 599 127 633 161
rect 599 59 633 93
rect 693 59 727 93
rect 787 127 821 161
rect 787 59 821 93
rect 881 59 915 93
rect 975 127 1009 161
rect 975 59 1009 93
rect 1069 59 1103 93
rect 1163 127 1197 161
rect 1163 59 1197 93
rect 1257 127 1291 161
rect 1351 59 1385 93
rect 1445 127 1479 161
rect 1539 59 1573 93
rect 1633 127 1667 161
rect 1727 59 1761 93
rect 1821 127 1855 161
rect 1915 59 1949 93
rect 2009 127 2043 161
rect 2103 59 2137 93
rect 2197 127 2231 161
rect 2291 127 2325 161
rect 2291 59 2325 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 505 451 539 485
rect 505 383 539 417
rect 505 315 539 349
rect 599 451 633 485
rect 599 383 633 417
rect 693 451 727 485
rect 693 383 727 417
rect 693 315 727 349
rect 787 451 821 485
rect 787 383 821 417
rect 881 451 915 485
rect 881 383 915 417
rect 881 315 915 349
rect 975 451 1009 485
rect 975 383 1009 417
rect 1069 451 1103 485
rect 1069 383 1103 417
rect 1069 315 1103 349
rect 1163 451 1197 485
rect 1163 383 1197 417
rect 1257 451 1291 485
rect 1257 383 1291 417
rect 1257 315 1291 349
rect 1351 451 1385 485
rect 1351 383 1385 417
rect 1445 451 1479 485
rect 1445 383 1479 417
rect 1445 315 1479 349
rect 1539 451 1573 485
rect 1539 383 1573 417
rect 1633 451 1667 485
rect 1633 383 1667 417
rect 1633 315 1667 349
rect 1727 451 1761 485
rect 1727 383 1761 417
rect 1821 451 1855 485
rect 1821 383 1855 417
rect 1821 315 1855 349
rect 1915 451 1949 485
rect 1915 383 1949 417
rect 2009 451 2043 485
rect 2009 383 2043 417
rect 2009 315 2043 349
rect 2103 451 2137 485
rect 2103 383 2137 417
rect 2197 451 2231 485
rect 2197 383 2231 417
rect 2197 315 2231 349
rect 2291 451 2325 485
rect 2291 383 2325 417
rect 2291 315 2325 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 1209 497 1245 523
rect 1303 497 1339 523
rect 1397 497 1433 523
rect 1491 497 1527 523
rect 1585 497 1621 523
rect 1679 497 1715 523
rect 1773 497 1809 523
rect 1867 497 1903 523
rect 1961 497 1997 523
rect 2055 497 2091 523
rect 2149 497 2185 523
rect 2243 497 2279 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 1209 282 1245 297
rect 1303 282 1339 297
rect 1397 282 1433 297
rect 1491 282 1527 297
rect 1585 282 1621 297
rect 1679 282 1715 297
rect 1773 282 1809 297
rect 1867 282 1903 297
rect 1961 282 1997 297
rect 2055 282 2091 297
rect 2149 282 2185 297
rect 2243 282 2279 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 831 265 871 282
rect 925 265 965 282
rect 1019 265 1059 282
rect 1113 265 1153 282
rect 67 249 1153 265
rect 67 215 83 249
rect 117 215 151 249
rect 185 215 219 249
rect 253 215 287 249
rect 321 215 355 249
rect 389 215 423 249
rect 457 215 491 249
rect 525 215 559 249
rect 593 215 627 249
rect 661 215 695 249
rect 729 215 763 249
rect 797 215 831 249
rect 865 215 899 249
rect 933 215 967 249
rect 1001 215 1035 249
rect 1069 215 1103 249
rect 1137 215 1153 249
rect 67 199 1153 215
rect 79 177 109 199
rect 183 177 213 199
rect 267 177 297 199
rect 371 177 401 199
rect 455 177 485 199
rect 559 177 589 199
rect 643 177 673 199
rect 747 177 777 199
rect 831 177 861 199
rect 935 177 965 199
rect 1019 177 1049 199
rect 1123 177 1153 199
rect 1207 265 1247 282
rect 1301 265 1341 282
rect 1395 265 1435 282
rect 1489 265 1529 282
rect 1583 265 1623 282
rect 1677 265 1717 282
rect 1771 265 1811 282
rect 1865 265 1905 282
rect 1959 265 1999 282
rect 2053 265 2093 282
rect 2147 265 2187 282
rect 2241 265 2281 282
rect 1207 249 2281 265
rect 1207 215 1341 249
rect 1375 215 1409 249
rect 1443 215 1477 249
rect 1511 215 1545 249
rect 1579 215 1613 249
rect 1647 215 1681 249
rect 1715 215 1749 249
rect 1783 215 1817 249
rect 1851 215 1885 249
rect 1919 215 1953 249
rect 1987 215 2021 249
rect 2055 215 2089 249
rect 2123 215 2281 249
rect 1207 199 2281 215
rect 1207 177 1237 199
rect 1301 177 1331 199
rect 1395 177 1425 199
rect 1499 177 1529 199
rect 1583 177 1613 199
rect 1687 177 1717 199
rect 1771 177 1801 199
rect 1865 177 1895 199
rect 1959 177 1989 199
rect 2063 177 2093 199
rect 2147 177 2177 199
rect 2251 177 2281 199
rect 79 21 109 47
rect 183 21 213 47
rect 267 21 297 47
rect 371 21 401 47
rect 455 21 485 47
rect 559 21 589 47
rect 643 21 673 47
rect 747 21 777 47
rect 831 21 861 47
rect 935 21 965 47
rect 1019 21 1049 47
rect 1123 21 1153 47
rect 1207 21 1237 47
rect 1301 21 1331 47
rect 1395 21 1425 47
rect 1499 21 1529 47
rect 1583 21 1613 47
rect 1687 21 1717 47
rect 1771 21 1801 47
rect 1865 21 1895 47
rect 1959 21 1989 47
rect 2063 21 2093 47
rect 2147 21 2177 47
rect 2251 21 2281 47
<< polycont >>
rect 83 215 117 249
rect 151 215 185 249
rect 219 215 253 249
rect 287 215 321 249
rect 355 215 389 249
rect 423 215 457 249
rect 491 215 525 249
rect 559 215 593 249
rect 627 215 661 249
rect 695 215 729 249
rect 763 215 797 249
rect 831 215 865 249
rect 899 215 933 249
rect 967 215 1001 249
rect 1035 215 1069 249
rect 1103 215 1137 249
rect 1341 215 1375 249
rect 1409 215 1443 249
rect 1477 215 1511 249
rect 1545 215 1579 249
rect 1613 215 1647 249
rect 1681 215 1715 249
rect 1749 215 1783 249
rect 1817 215 1851 249
rect 1885 215 1919 249
rect 1953 215 1987 249
rect 2021 215 2055 249
rect 2089 215 2123 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 25 485 79 527
rect 25 451 35 485
rect 69 451 79 485
rect 25 417 79 451
rect 25 383 35 417
rect 69 383 79 417
rect 25 349 79 383
rect 25 315 35 349
rect 69 315 79 349
rect 25 299 79 315
rect 113 485 179 493
rect 113 451 129 485
rect 163 451 179 485
rect 113 417 179 451
rect 113 383 129 417
rect 163 383 179 417
rect 113 349 179 383
rect 213 485 267 527
rect 213 451 223 485
rect 257 451 267 485
rect 213 417 267 451
rect 213 383 223 417
rect 257 383 267 417
rect 213 367 267 383
rect 301 485 367 493
rect 301 451 317 485
rect 351 451 367 485
rect 301 417 367 451
rect 301 383 317 417
rect 351 383 367 417
rect 113 315 129 349
rect 163 333 179 349
rect 301 349 367 383
rect 401 485 455 527
rect 401 451 411 485
rect 445 451 455 485
rect 401 417 455 451
rect 401 383 411 417
rect 445 383 455 417
rect 401 367 455 383
rect 489 485 555 493
rect 489 451 505 485
rect 539 451 555 485
rect 489 417 555 451
rect 489 383 505 417
rect 539 383 555 417
rect 301 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 489 349 555 383
rect 589 485 643 527
rect 589 451 599 485
rect 633 451 643 485
rect 589 417 643 451
rect 589 383 599 417
rect 633 383 643 417
rect 589 367 643 383
rect 677 485 743 493
rect 677 451 693 485
rect 727 451 743 485
rect 677 417 743 451
rect 677 383 693 417
rect 727 383 743 417
rect 489 333 505 349
rect 351 315 505 333
rect 539 333 555 349
rect 677 349 743 383
rect 777 485 831 527
rect 777 451 787 485
rect 821 451 831 485
rect 777 417 831 451
rect 777 383 787 417
rect 821 383 831 417
rect 777 367 831 383
rect 865 485 931 493
rect 865 451 881 485
rect 915 451 931 485
rect 865 417 931 451
rect 865 383 881 417
rect 915 383 931 417
rect 677 333 693 349
rect 539 315 693 333
rect 727 333 743 349
rect 865 349 931 383
rect 965 485 1019 527
rect 965 451 975 485
rect 1009 451 1019 485
rect 965 417 1019 451
rect 965 383 975 417
rect 1009 383 1019 417
rect 965 367 1019 383
rect 1053 485 1119 493
rect 1053 451 1069 485
rect 1103 451 1119 485
rect 1053 417 1119 451
rect 1053 383 1069 417
rect 1103 383 1119 417
rect 865 333 881 349
rect 727 315 881 333
rect 915 333 931 349
rect 1053 349 1119 383
rect 1153 485 1207 527
rect 1153 451 1163 485
rect 1197 451 1207 485
rect 1153 417 1207 451
rect 1153 383 1163 417
rect 1197 383 1207 417
rect 1153 367 1207 383
rect 1241 485 1307 493
rect 1241 451 1257 485
rect 1291 451 1307 485
rect 1241 417 1307 451
rect 1241 383 1257 417
rect 1291 383 1307 417
rect 1053 333 1069 349
rect 915 315 1069 333
rect 1103 333 1119 349
rect 1241 349 1307 383
rect 1341 485 1395 527
rect 1341 451 1351 485
rect 1385 451 1395 485
rect 1341 417 1395 451
rect 1341 383 1351 417
rect 1385 383 1395 417
rect 1341 367 1395 383
rect 1429 485 1495 493
rect 1429 451 1445 485
rect 1479 451 1495 485
rect 1429 417 1495 451
rect 1429 383 1445 417
rect 1479 383 1495 417
rect 1241 333 1257 349
rect 1103 315 1257 333
rect 1291 333 1307 349
rect 1429 349 1495 383
rect 1529 485 1583 527
rect 1529 451 1539 485
rect 1573 451 1583 485
rect 1529 417 1583 451
rect 1529 383 1539 417
rect 1573 383 1583 417
rect 1529 367 1583 383
rect 1617 485 1683 493
rect 1617 451 1633 485
rect 1667 451 1683 485
rect 1617 417 1683 451
rect 1617 383 1633 417
rect 1667 383 1683 417
rect 1429 333 1445 349
rect 1291 315 1445 333
rect 1479 333 1495 349
rect 1617 349 1683 383
rect 1717 485 1771 527
rect 1717 451 1727 485
rect 1761 451 1771 485
rect 1717 417 1771 451
rect 1717 383 1727 417
rect 1761 383 1771 417
rect 1717 367 1771 383
rect 1805 485 1871 493
rect 1805 451 1821 485
rect 1855 451 1871 485
rect 1805 417 1871 451
rect 1805 383 1821 417
rect 1855 383 1871 417
rect 1617 333 1633 349
rect 1479 315 1633 333
rect 1667 333 1683 349
rect 1805 349 1871 383
rect 1905 485 1959 527
rect 1905 451 1915 485
rect 1949 451 1959 485
rect 1905 417 1959 451
rect 1905 383 1915 417
rect 1949 383 1959 417
rect 1905 367 1959 383
rect 1993 485 2059 493
rect 1993 451 2009 485
rect 2043 451 2059 485
rect 1993 417 2059 451
rect 1993 383 2009 417
rect 2043 383 2059 417
rect 1805 333 1821 349
rect 1667 315 1821 333
rect 1855 333 1871 349
rect 1993 349 2059 383
rect 2093 485 2147 527
rect 2093 451 2103 485
rect 2137 451 2147 485
rect 2093 417 2147 451
rect 2093 383 2103 417
rect 2137 383 2147 417
rect 2093 367 2147 383
rect 2181 485 2247 493
rect 2181 451 2197 485
rect 2231 451 2247 485
rect 2181 417 2247 451
rect 2181 383 2197 417
rect 2231 383 2247 417
rect 1993 333 2009 349
rect 1855 315 2009 333
rect 2043 333 2059 349
rect 2181 349 2247 383
rect 2181 333 2197 349
rect 2043 315 2197 333
rect 2231 315 2247 349
rect 113 299 2247 315
rect 2281 485 2335 527
rect 2281 451 2291 485
rect 2325 451 2335 485
rect 2281 417 2335 451
rect 2281 383 2291 417
rect 2325 383 2335 417
rect 2281 349 2335 383
rect 2281 315 2291 349
rect 2325 315 2335 349
rect 2281 299 2335 315
rect 67 249 1153 265
rect 67 215 83 249
rect 117 215 151 249
rect 185 215 219 249
rect 253 215 287 249
rect 321 215 355 249
rect 389 215 423 249
rect 457 215 491 249
rect 525 215 559 249
rect 593 215 627 249
rect 661 215 695 249
rect 729 215 763 249
rect 797 215 831 249
rect 865 215 899 249
rect 933 215 967 249
rect 1001 215 1035 249
rect 1069 215 1103 249
rect 1137 215 1153 249
rect 67 211 1153 215
rect 1209 211 1291 299
rect 2193 265 2247 299
rect 1325 249 2139 265
rect 1325 215 1341 249
rect 1375 215 1409 249
rect 1443 215 1477 249
rect 1511 215 1545 249
rect 1579 215 1613 249
rect 1647 215 1681 249
rect 1715 215 1749 249
rect 1783 215 1817 249
rect 1851 215 1885 249
rect 1919 215 1953 249
rect 1987 215 2021 249
rect 2055 215 2089 249
rect 2123 215 2139 249
rect 1325 211 2139 215
rect 2193 211 2287 265
rect 1231 177 1291 211
rect 2193 177 2247 211
rect 18 161 1197 177
rect 18 127 35 161
rect 69 143 223 161
rect 69 127 85 143
rect 18 93 85 127
rect 207 127 223 143
rect 257 143 411 161
rect 257 127 273 143
rect 18 59 35 93
rect 69 59 85 93
rect 18 51 85 59
rect 119 93 173 109
rect 119 59 129 93
rect 163 59 173 93
rect 119 17 173 59
rect 207 93 273 127
rect 395 127 411 143
rect 445 143 599 161
rect 445 127 461 143
rect 207 59 223 93
rect 257 59 273 93
rect 207 51 273 59
rect 307 93 361 109
rect 307 59 317 93
rect 351 59 361 93
rect 307 17 361 59
rect 395 93 461 127
rect 583 127 599 143
rect 633 143 787 161
rect 633 127 649 143
rect 395 59 411 93
rect 445 59 461 93
rect 395 51 461 59
rect 495 93 549 109
rect 495 59 505 93
rect 539 59 549 93
rect 495 17 549 59
rect 583 93 649 127
rect 771 127 787 143
rect 821 143 975 161
rect 821 127 837 143
rect 583 59 599 93
rect 633 59 649 93
rect 583 51 649 59
rect 683 93 737 109
rect 683 59 693 93
rect 727 59 737 93
rect 683 17 737 59
rect 771 93 837 127
rect 959 127 975 143
rect 1009 143 1163 161
rect 1009 127 1025 143
rect 771 59 787 93
rect 821 59 837 93
rect 771 51 837 59
rect 871 93 925 109
rect 871 59 881 93
rect 915 59 925 93
rect 871 17 925 59
rect 959 93 1025 127
rect 1147 127 1163 143
rect 1231 161 2247 177
rect 1231 127 1257 161
rect 1291 127 1445 161
rect 1479 127 1633 161
rect 1667 127 1821 161
rect 1855 127 2009 161
rect 2043 127 2197 161
rect 2231 127 2247 161
rect 2291 161 2341 177
rect 2325 127 2341 161
rect 959 59 975 93
rect 1009 59 1025 93
rect 959 51 1025 59
rect 1059 93 1113 109
rect 1059 59 1069 93
rect 1103 59 1113 93
rect 1059 17 1113 59
rect 1147 93 1197 127
rect 2291 93 2341 127
rect 1147 59 1163 93
rect 1197 59 1351 93
rect 1385 59 1539 93
rect 1573 59 1727 93
rect 1761 59 1915 93
rect 1949 59 2103 93
rect 2137 59 2291 93
rect 2325 59 2341 93
rect 1147 51 2341 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< labels >>
flabel locali s 1225 221 1259 255 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 1777 221 1811 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2_12
<< properties >>
string FIXED_BBOX 0 0 2392 544
string GDS_END 308474
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 291458
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
