magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 2890 582
<< pwell >>
rect 1538 157 1939 201
rect 2528 157 2835 203
rect 1 21 2835 157
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 131
rect 171 47 201 131
rect 265 47 295 131
rect 349 47 379 131
rect 563 47 593 131
rect 761 47 791 131
rect 855 47 885 131
rect 1053 47 1083 131
rect 1147 47 1177 131
rect 1229 47 1259 131
rect 1437 47 1467 131
rect 1519 47 1549 131
rect 1624 47 1654 175
rect 1813 47 1843 175
rect 1965 47 1995 131
rect 2037 47 2067 131
rect 2163 47 2193 131
rect 2287 47 2317 131
rect 2509 47 2539 131
rect 2614 47 2644 177
rect 2708 47 2738 177
<< scpmoshvt >>
rect 81 369 117 497
rect 175 369 211 497
rect 257 369 293 497
rect 351 369 387 497
rect 549 369 585 497
rect 747 369 783 497
rect 841 369 877 497
rect 1039 413 1075 497
rect 1133 413 1169 497
rect 1245 413 1281 497
rect 1383 413 1419 497
rect 1501 413 1537 497
rect 1627 329 1663 497
rect 1709 329 1745 497
rect 1855 413 1891 497
rect 1953 413 1989 497
rect 2095 413 2131 497
rect 2303 413 2339 497
rect 2501 369 2537 497
rect 2606 297 2642 497
rect 2700 297 2736 497
<< ndiff >>
rect 1564 131 1624 175
rect 27 103 89 131
rect 27 69 35 103
rect 69 69 89 103
rect 27 47 89 69
rect 119 47 171 131
rect 201 93 265 131
rect 201 59 211 93
rect 245 59 265 93
rect 201 47 265 59
rect 295 47 349 131
rect 379 93 447 131
rect 379 59 405 93
rect 439 59 447 93
rect 379 47 447 59
rect 501 105 563 131
rect 501 71 509 105
rect 543 71 563 105
rect 501 47 563 71
rect 593 93 645 131
rect 593 59 603 93
rect 637 59 645 93
rect 593 47 645 59
rect 699 105 761 131
rect 699 71 707 105
rect 741 71 761 105
rect 699 47 761 71
rect 791 89 855 131
rect 791 55 801 89
rect 835 55 855 89
rect 791 47 855 55
rect 885 101 937 131
rect 885 67 895 101
rect 929 67 937 101
rect 885 47 937 67
rect 991 101 1053 131
rect 991 67 999 101
rect 1033 67 1053 101
rect 991 47 1053 67
rect 1083 101 1147 131
rect 1083 67 1093 101
rect 1127 67 1147 101
rect 1083 47 1147 67
rect 1177 47 1229 131
rect 1259 93 1311 131
rect 1259 59 1269 93
rect 1303 59 1311 93
rect 1259 47 1311 59
rect 1365 119 1437 131
rect 1365 85 1373 119
rect 1407 85 1437 119
rect 1365 47 1437 85
rect 1467 47 1519 131
rect 1549 89 1624 131
rect 1549 55 1561 89
rect 1595 55 1624 89
rect 1549 47 1624 55
rect 1654 47 1813 175
rect 1843 131 1913 175
rect 2554 131 2614 177
rect 1843 89 1965 131
rect 1843 55 1869 89
rect 1903 55 1965 89
rect 1843 47 1965 55
rect 1995 47 2037 131
rect 2067 47 2163 131
rect 2193 89 2287 131
rect 2193 55 2233 89
rect 2267 55 2287 89
rect 2193 47 2287 55
rect 2317 101 2393 131
rect 2317 67 2351 101
rect 2385 67 2393 101
rect 2317 47 2393 67
rect 2447 102 2509 131
rect 2447 68 2455 102
rect 2489 68 2509 102
rect 2447 47 2509 68
rect 2539 89 2614 131
rect 2539 55 2554 89
rect 2588 55 2614 89
rect 2539 47 2614 55
rect 2644 105 2708 177
rect 2644 71 2654 105
rect 2688 71 2708 105
rect 2644 47 2708 71
rect 2738 161 2809 177
rect 2738 127 2765 161
rect 2799 127 2809 161
rect 2738 93 2809 127
rect 2738 59 2765 93
rect 2799 59 2809 93
rect 2738 47 2809 59
<< pdiff >>
rect 27 431 81 497
rect 27 397 35 431
rect 69 397 81 431
rect 27 369 81 397
rect 117 489 175 497
rect 117 455 129 489
rect 163 455 175 489
rect 117 369 175 455
rect 211 369 257 497
rect 293 411 351 497
rect 293 377 305 411
rect 339 377 351 411
rect 293 369 351 377
rect 387 485 441 497
rect 387 451 399 485
rect 433 451 441 485
rect 387 369 441 451
rect 495 415 549 497
rect 495 381 503 415
rect 537 381 549 415
rect 495 369 549 381
rect 585 485 639 497
rect 585 451 597 485
rect 631 451 639 485
rect 585 369 639 451
rect 693 449 747 497
rect 693 415 701 449
rect 735 415 747 449
rect 693 369 747 415
rect 783 489 841 497
rect 783 455 795 489
rect 829 455 841 489
rect 783 369 841 455
rect 877 477 931 497
rect 877 443 889 477
rect 923 443 931 477
rect 877 369 931 443
rect 985 477 1039 497
rect 985 443 993 477
rect 1027 443 1039 477
rect 985 413 1039 443
rect 1075 477 1133 497
rect 1075 443 1087 477
rect 1121 443 1133 477
rect 1075 413 1133 443
rect 1169 413 1245 497
rect 1281 489 1383 497
rect 1281 455 1305 489
rect 1339 455 1383 489
rect 1281 413 1383 455
rect 1419 474 1501 497
rect 1419 440 1436 474
rect 1470 440 1501 474
rect 1419 413 1501 440
rect 1537 489 1627 497
rect 1537 455 1558 489
rect 1592 455 1627 489
rect 1537 413 1627 455
rect 1575 329 1627 413
rect 1663 329 1709 497
rect 1745 475 1855 497
rect 1745 441 1787 475
rect 1821 441 1855 475
rect 1745 413 1855 441
rect 1891 413 1953 497
rect 1989 489 2095 497
rect 1989 455 2028 489
rect 2062 455 2095 489
rect 1989 413 2095 455
rect 2131 474 2195 497
rect 2131 440 2143 474
rect 2177 440 2195 474
rect 2131 413 2195 440
rect 2249 485 2303 497
rect 2249 451 2257 485
rect 2291 451 2303 485
rect 2249 413 2303 451
rect 2339 474 2393 497
rect 2339 440 2351 474
rect 2385 440 2393 474
rect 2339 413 2393 440
rect 2447 483 2501 497
rect 2447 449 2455 483
rect 2489 449 2501 483
rect 2447 415 2501 449
rect 1745 329 1797 413
rect 2447 381 2455 415
rect 2489 381 2501 415
rect 2447 369 2501 381
rect 2537 489 2606 497
rect 2537 455 2554 489
rect 2588 455 2606 489
rect 2537 421 2606 455
rect 2537 387 2554 421
rect 2588 387 2606 421
rect 2537 369 2606 387
rect 2554 297 2606 369
rect 2642 474 2700 497
rect 2642 440 2654 474
rect 2688 440 2700 474
rect 2642 297 2700 440
rect 2736 485 2809 497
rect 2736 451 2765 485
rect 2799 451 2809 485
rect 2736 417 2809 451
rect 2736 383 2765 417
rect 2799 383 2809 417
rect 2736 349 2809 383
rect 2736 315 2765 349
rect 2799 315 2809 349
rect 2736 297 2809 315
<< ndiffc >>
rect 35 69 69 103
rect 211 59 245 93
rect 405 59 439 93
rect 509 71 543 105
rect 603 59 637 93
rect 707 71 741 105
rect 801 55 835 89
rect 895 67 929 101
rect 999 67 1033 101
rect 1093 67 1127 101
rect 1269 59 1303 93
rect 1373 85 1407 119
rect 1561 55 1595 89
rect 1869 55 1903 89
rect 2233 55 2267 89
rect 2351 67 2385 101
rect 2455 68 2489 102
rect 2554 55 2588 89
rect 2654 71 2688 105
rect 2765 127 2799 161
rect 2765 59 2799 93
<< pdiffc >>
rect 35 397 69 431
rect 129 455 163 489
rect 305 377 339 411
rect 399 451 433 485
rect 503 381 537 415
rect 597 451 631 485
rect 701 415 735 449
rect 795 455 829 489
rect 889 443 923 477
rect 993 443 1027 477
rect 1087 443 1121 477
rect 1305 455 1339 489
rect 1436 440 1470 474
rect 1558 455 1592 489
rect 1787 441 1821 475
rect 2028 455 2062 489
rect 2143 440 2177 474
rect 2257 451 2291 485
rect 2351 440 2385 474
rect 2455 449 2489 483
rect 2455 381 2489 415
rect 2554 455 2588 489
rect 2554 387 2588 421
rect 2654 440 2688 474
rect 2765 451 2799 485
rect 2765 383 2799 417
rect 2765 315 2799 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 257 497 293 523
rect 351 497 387 523
rect 549 497 585 523
rect 747 497 783 523
rect 841 497 877 523
rect 1039 497 1075 523
rect 1133 497 1169 523
rect 1245 497 1281 523
rect 1383 497 1419 523
rect 1501 497 1537 523
rect 1627 497 1663 523
rect 1709 497 1745 523
rect 1855 497 1891 523
rect 1953 497 1989 523
rect 2095 497 2131 523
rect 2303 497 2339 523
rect 2501 497 2537 523
rect 2606 497 2642 523
rect 2700 497 2736 523
rect 1039 398 1075 413
rect 1133 398 1169 413
rect 1245 398 1281 413
rect 1383 398 1419 413
rect 1501 398 1537 413
rect 81 354 117 369
rect 175 354 211 369
rect 257 354 293 369
rect 351 354 387 369
rect 549 354 585 369
rect 747 354 783 369
rect 841 354 877 369
rect 978 368 1077 398
rect 1131 381 1171 398
rect 1243 381 1283 398
rect 48 324 119 354
rect 48 265 78 324
rect 173 283 213 354
rect 21 249 78 265
rect 21 215 34 249
rect 68 215 78 249
rect 130 267 213 283
rect 130 233 140 267
rect 174 253 213 267
rect 174 233 201 253
rect 130 217 201 233
rect 255 219 295 354
rect 349 265 389 354
rect 547 265 587 354
rect 733 324 785 354
rect 733 284 763 324
rect 839 284 879 354
rect 978 284 1008 368
rect 1119 365 1183 381
rect 1119 331 1129 365
rect 1163 331 1183 365
rect 1119 315 1183 331
rect 1243 365 1329 381
rect 1243 331 1285 365
rect 1319 331 1329 365
rect 1243 315 1329 331
rect 709 268 763 284
rect 349 249 478 265
rect 21 199 78 215
rect 48 176 78 199
rect 48 146 119 176
rect 89 131 119 146
rect 171 131 201 217
rect 243 203 307 219
rect 243 169 253 203
rect 287 169 307 203
rect 243 153 307 169
rect 349 215 413 249
rect 447 215 478 249
rect 349 199 478 215
rect 520 249 593 265
rect 520 215 530 249
rect 564 215 593 249
rect 709 234 719 268
rect 753 234 763 268
rect 709 218 763 234
rect 815 268 879 284
rect 815 234 825 268
rect 859 234 879 268
rect 815 218 879 234
rect 924 268 1008 284
rect 924 234 934 268
rect 968 248 1008 268
rect 968 234 1177 248
rect 924 218 1177 234
rect 520 199 593 215
rect 265 131 295 153
rect 349 131 379 199
rect 563 131 593 199
rect 733 176 763 218
rect 842 176 879 218
rect 733 146 791 176
rect 842 146 1083 176
rect 761 131 791 146
rect 855 131 885 146
rect 1053 131 1083 146
rect 1147 131 1177 218
rect 1243 213 1283 315
rect 1381 273 1421 398
rect 1499 369 1539 398
rect 1473 353 1539 369
rect 1473 319 1483 353
rect 1517 319 1539 353
rect 1855 398 1891 413
rect 1953 398 1989 413
rect 2095 398 2131 413
rect 2303 398 2339 413
rect 1853 381 1893 398
rect 1835 365 1909 381
rect 1835 345 1855 365
rect 1813 331 1855 345
rect 1889 331 1909 365
rect 1473 303 1539 319
rect 1627 314 1663 329
rect 1709 314 1745 329
rect 1813 315 1909 331
rect 1951 325 1991 398
rect 2093 397 2133 398
rect 2093 367 2193 397
rect 2119 343 2193 367
rect 2301 365 2341 398
rect 1345 263 1421 273
rect 1345 229 1361 263
rect 1395 229 1421 263
rect 1499 273 1539 303
rect 1499 243 1549 273
rect 1625 265 1665 314
rect 1345 219 1421 229
rect 1229 203 1295 213
rect 1229 169 1245 203
rect 1279 169 1295 203
rect 1229 159 1295 169
rect 1381 176 1421 219
rect 1229 131 1259 159
rect 1381 146 1467 176
rect 1437 131 1467 146
rect 1519 131 1549 243
rect 1591 249 1665 265
rect 1591 215 1601 249
rect 1635 215 1665 249
rect 1591 199 1665 215
rect 1707 265 1747 314
rect 1707 249 1771 265
rect 1707 215 1717 249
rect 1751 215 1771 249
rect 1707 199 1771 215
rect 1624 175 1654 199
rect 1813 175 1843 315
rect 1951 295 2077 325
rect 1931 235 1995 251
rect 1931 201 1941 235
rect 1975 201 1995 235
rect 1931 185 1995 201
rect 1965 131 1995 185
rect 2037 237 2077 295
rect 2119 309 2139 343
rect 2173 309 2193 343
rect 2241 355 2341 365
rect 2241 321 2257 355
rect 2291 321 2341 355
rect 2501 354 2537 369
rect 2241 311 2341 321
rect 2119 293 2193 309
rect 2037 221 2101 237
rect 2037 187 2047 221
rect 2081 187 2101 221
rect 2037 171 2101 187
rect 2037 131 2067 171
rect 2163 131 2193 293
rect 2253 271 2341 311
rect 2499 271 2539 354
rect 2606 282 2642 297
rect 2700 282 2736 297
rect 2253 241 2539 271
rect 2604 265 2644 282
rect 2698 265 2738 282
rect 2253 203 2317 241
rect 2253 169 2263 203
rect 2297 169 2317 203
rect 2253 153 2317 169
rect 2287 131 2317 153
rect 2509 131 2539 241
rect 2581 249 2738 265
rect 2581 215 2591 249
rect 2625 215 2738 249
rect 2581 199 2738 215
rect 2614 177 2644 199
rect 2708 177 2738 199
rect 89 21 119 47
rect 171 21 201 47
rect 265 21 295 47
rect 349 21 379 47
rect 563 21 593 47
rect 761 21 791 47
rect 855 21 885 47
rect 1053 21 1083 47
rect 1147 21 1177 47
rect 1229 21 1259 47
rect 1437 21 1467 47
rect 1519 21 1549 47
rect 1624 21 1654 47
rect 1813 21 1843 47
rect 1965 21 1995 47
rect 2037 21 2067 47
rect 2163 21 2193 47
rect 2287 21 2317 47
rect 2509 21 2539 47
rect 2614 21 2644 47
rect 2708 21 2738 47
<< polycont >>
rect 34 215 68 249
rect 140 233 174 267
rect 1129 331 1163 365
rect 1285 331 1319 365
rect 253 169 287 203
rect 413 215 447 249
rect 530 215 564 249
rect 719 234 753 268
rect 825 234 859 268
rect 934 234 968 268
rect 1483 319 1517 353
rect 1855 331 1889 365
rect 1361 229 1395 263
rect 1245 169 1279 203
rect 1601 215 1635 249
rect 1717 215 1751 249
rect 1941 201 1975 235
rect 2139 309 2173 343
rect 2257 321 2291 355
rect 2047 187 2081 221
rect 2263 169 2297 203
rect 2591 215 2625 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 17 431 69 493
rect 103 489 167 527
rect 103 455 129 489
rect 163 455 167 489
rect 103 439 167 455
rect 211 485 449 493
rect 211 451 399 485
rect 433 451 449 485
rect 17 397 35 431
rect 211 405 245 451
rect 494 417 544 493
rect 588 485 647 527
rect 588 451 597 485
rect 631 451 647 485
rect 769 489 845 527
rect 588 428 647 451
rect 701 449 735 465
rect 769 455 795 489
rect 829 455 845 489
rect 889 477 958 493
rect 69 397 245 405
rect 17 369 245 397
rect 279 411 369 417
rect 279 377 305 411
rect 339 377 369 411
rect 279 369 369 377
rect 17 249 68 335
rect 17 215 34 249
rect 17 153 68 215
rect 108 267 174 335
rect 108 255 140 267
rect 108 221 128 255
rect 162 221 174 233
rect 108 153 174 221
rect 208 203 297 335
rect 208 169 253 203
rect 287 169 297 203
rect 208 153 297 169
rect 331 323 369 369
rect 331 289 335 323
rect 331 119 369 289
rect 413 415 544 417
rect 413 381 503 415
rect 537 381 544 415
rect 413 354 544 381
rect 923 443 958 477
rect 889 427 958 443
rect 701 400 735 415
rect 701 391 859 400
rect 701 366 825 391
rect 807 357 825 366
rect 413 249 480 354
rect 447 215 480 249
rect 514 255 590 320
rect 514 221 529 255
rect 563 249 590 255
rect 514 215 530 221
rect 564 215 590 249
rect 631 268 763 330
rect 631 234 719 268
rect 753 234 763 268
rect 413 181 480 215
rect 631 211 763 234
rect 807 268 859 357
rect 807 234 825 268
rect 413 143 544 181
rect 807 177 859 234
rect 17 103 150 119
rect 17 69 35 103
rect 69 69 150 103
rect 17 17 150 69
rect 184 93 369 119
rect 184 59 211 93
rect 245 59 369 93
rect 184 51 369 59
rect 405 93 458 109
rect 439 59 458 93
rect 405 17 458 59
rect 492 105 544 143
rect 704 143 859 177
rect 895 284 958 427
rect 993 477 1036 493
rect 1027 443 1036 477
rect 993 323 1036 443
rect 1087 477 1241 493
rect 1121 443 1241 477
rect 1289 489 1366 527
rect 1289 455 1305 489
rect 1339 455 1366 489
rect 1431 474 1484 490
rect 1087 427 1241 443
rect 993 318 1002 323
rect 1155 365 1173 391
rect 1121 331 1129 357
rect 1163 331 1173 365
rect 1121 315 1173 331
rect 895 268 968 284
rect 895 254 934 268
rect 895 220 927 254
rect 961 220 968 234
rect 895 217 968 220
rect 492 71 509 105
rect 543 71 544 105
rect 492 51 544 71
rect 588 93 670 111
rect 588 59 603 93
rect 637 59 670 93
rect 588 17 670 59
rect 704 105 741 143
rect 704 71 707 105
rect 704 51 741 71
rect 785 89 851 109
rect 785 55 801 89
rect 835 55 851 89
rect 785 17 851 55
rect 895 101 937 217
rect 1002 156 1036 289
rect 1207 279 1241 427
rect 1431 440 1436 474
rect 1470 440 1484 474
rect 1431 421 1484 440
rect 1542 489 1753 527
rect 1542 455 1558 489
rect 1592 455 1753 489
rect 1542 425 1753 455
rect 1787 475 1968 492
rect 1821 441 1968 475
rect 2012 489 2088 527
rect 2012 455 2028 489
rect 2062 455 2088 489
rect 2012 447 2088 455
rect 2122 474 2203 490
rect 1787 425 1968 441
rect 1285 387 1484 421
rect 1934 413 1968 425
rect 2122 440 2143 474
rect 2177 440 2203 474
rect 2241 485 2317 527
rect 2241 451 2257 485
rect 2291 451 2317 485
rect 2241 447 2317 451
rect 2351 474 2403 493
rect 2122 413 2203 440
rect 2385 440 2403 474
rect 1285 365 1319 387
rect 1577 357 1642 391
rect 1676 357 1777 391
rect 1285 315 1319 331
rect 1438 319 1483 353
rect 1517 323 1543 353
rect 1577 334 1777 357
rect 1438 289 1487 319
rect 1521 289 1543 323
rect 929 67 937 101
rect 895 51 937 67
rect 971 101 1036 156
rect 971 67 999 101
rect 1033 67 1036 101
rect 971 51 1036 67
rect 1093 263 1395 279
rect 1093 245 1361 263
rect 1093 101 1178 245
rect 1601 255 1683 265
rect 1395 249 1683 255
rect 1395 229 1601 249
rect 1361 215 1601 229
rect 1635 215 1683 249
rect 1219 169 1245 203
rect 1279 169 1295 203
rect 1361 195 1683 215
rect 1717 249 1777 334
rect 1751 215 1777 249
rect 1835 365 1900 381
rect 1934 379 2317 413
rect 1835 331 1855 365
rect 1889 331 1900 365
rect 2241 355 2317 379
rect 1835 255 1900 331
rect 1946 343 2199 345
rect 1946 323 2139 343
rect 1946 289 1958 323
rect 1992 309 2139 323
rect 2173 309 2199 343
rect 2241 321 2257 355
rect 2291 321 2317 355
rect 1992 289 2007 309
rect 1946 285 2007 289
rect 2351 273 2403 440
rect 1835 221 1856 255
rect 1890 221 1900 255
rect 1835 215 1900 221
rect 1934 235 2001 251
rect 1219 161 1295 169
rect 1717 181 1777 215
rect 1934 201 1941 235
rect 1975 201 2001 235
rect 1934 181 2001 201
rect 1219 127 1407 161
rect 1127 67 1178 101
rect 1357 119 1407 127
rect 1093 51 1178 67
rect 1212 59 1269 93
rect 1303 59 1319 93
rect 1212 17 1319 59
rect 1357 85 1373 119
rect 1357 51 1407 85
rect 1451 89 1683 161
rect 1717 144 2001 181
rect 2044 239 2403 273
rect 2044 221 2096 239
rect 2044 187 2047 221
rect 2081 187 2096 221
rect 2044 171 2096 187
rect 2142 169 2263 203
rect 2297 169 2323 203
rect 2142 157 2323 169
rect 2142 109 2182 157
rect 2357 117 2403 239
rect 1451 55 1561 89
rect 1595 55 1683 89
rect 1853 89 2182 109
rect 1853 55 1869 89
rect 1903 55 2182 89
rect 2233 89 2283 109
rect 2267 55 2283 89
rect 1451 17 1683 55
rect 2233 17 2283 55
rect 2335 101 2403 117
rect 2335 67 2351 101
rect 2385 67 2403 101
rect 2335 51 2403 67
rect 2437 483 2505 493
rect 2437 449 2455 483
rect 2489 449 2505 483
rect 2437 415 2505 449
rect 2437 381 2455 415
rect 2489 381 2505 415
rect 2437 265 2505 381
rect 2553 489 2604 527
rect 2553 455 2554 489
rect 2588 455 2604 489
rect 2553 421 2604 455
rect 2553 387 2554 421
rect 2588 387 2604 421
rect 2553 369 2604 387
rect 2649 474 2731 490
rect 2649 440 2654 474
rect 2688 440 2731 474
rect 2649 299 2731 440
rect 2765 485 2799 527
rect 2765 417 2799 451
rect 2765 349 2799 383
rect 2765 299 2799 315
rect 2437 249 2625 265
rect 2437 215 2591 249
rect 2437 199 2625 215
rect 2437 102 2489 199
rect 2670 165 2731 299
rect 2437 68 2455 102
rect 2437 51 2489 68
rect 2523 89 2604 110
rect 2523 55 2554 89
rect 2588 55 2604 89
rect 2649 105 2731 165
rect 2649 71 2654 105
rect 2688 71 2731 105
rect 2649 55 2731 71
rect 2765 161 2799 177
rect 2765 93 2799 127
rect 2523 17 2604 55
rect 2765 17 2799 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 128 233 140 255
rect 140 233 162 255
rect 128 221 162 233
rect 335 289 369 323
rect 825 357 859 391
rect 529 249 563 255
rect 529 221 530 249
rect 530 221 563 249
rect 1002 289 1036 323
rect 1121 365 1155 391
rect 1121 357 1129 365
rect 1129 357 1155 365
rect 927 234 934 254
rect 934 234 961 254
rect 927 220 961 234
rect 1642 357 1676 391
rect 1487 319 1517 323
rect 1517 319 1521 323
rect 1487 289 1521 319
rect 1958 289 1992 323
rect 1856 221 1890 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
<< metal1 >>
rect 0 561 2852 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 0 496 2852 527
rect 813 391 881 397
rect 813 357 825 391
rect 859 388 881 391
rect 1109 391 1177 397
rect 1109 388 1121 391
rect 859 360 1121 388
rect 859 357 881 360
rect 813 351 881 357
rect 1109 357 1121 360
rect 1155 388 1177 391
rect 1630 391 1698 397
rect 1630 388 1642 391
rect 1155 360 1642 388
rect 1155 357 1177 360
rect 1109 351 1177 357
rect 1630 357 1642 360
rect 1676 357 1698 391
rect 1630 351 1698 357
rect 323 323 391 329
rect 323 289 335 323
rect 369 320 391 323
rect 990 323 1048 329
rect 990 320 1002 323
rect 369 292 1002 320
rect 369 289 391 292
rect 323 283 391 289
rect 990 289 1002 292
rect 1036 289 1048 323
rect 990 283 1048 289
rect 1475 323 1543 329
rect 1475 289 1487 323
rect 1521 320 1543 323
rect 1946 323 2014 329
rect 1946 320 1958 323
rect 1521 292 1958 320
rect 1521 289 1543 292
rect 1475 283 1543 289
rect 1946 289 1958 292
rect 1992 289 2014 323
rect 1946 283 2014 289
rect 116 255 174 261
rect 116 221 128 255
rect 162 252 174 255
rect 517 255 575 261
rect 517 252 529 255
rect 162 224 529 252
rect 162 221 174 224
rect 116 215 174 221
rect 517 221 529 224
rect 563 221 575 255
rect 517 215 575 221
rect 915 254 973 260
rect 915 220 927 254
rect 961 252 973 254
rect 1834 255 1912 261
rect 1834 252 1856 255
rect 961 224 1856 252
rect 961 220 973 224
rect 915 214 973 220
rect 1834 221 1856 224
rect 1890 221 1912 255
rect 1834 215 1912 221
rect 0 17 2852 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
rect 0 -48 2852 -17
<< labels >>
flabel locali s 2673 289 2707 323 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2673 85 2707 119 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2673 153 2707 187 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2673 221 2707 255 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2673 425 2707 459 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2673 357 2707 391 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 SCD
port 3 nsew signal input
flabel locali s 213 289 247 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 SCD
port 3 nsew signal input
flabel locali s 213 153 247 187 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew signal input
flabel metal1 s 1501 289 1535 323 0 FreeSans 200 0 0 0 SET_B
port 5 nsew signal input
flabel metal1 s 121 221 155 255 0 FreeSans 200 0 0 0 SCE
port 4 nsew signal input
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel comment s 2309 287 2309 287 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfstp_4
flabel comment s 1263 286 1263 286 0 FreeSans 200 0 0 0 no_jumper_check
<< properties >>
string FIXED_BBOX 0 0 2852 544
string GDS_END 2575374
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 2555046
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
