magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1909 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 287 47 317 177
rect 381 47 411 177
rect 475 47 505 177
rect 569 47 599 177
rect 663 47 693 177
rect 757 47 787 177
rect 851 47 881 177
rect 945 47 975 177
rect 1143 47 1173 177
rect 1237 47 1267 177
rect 1331 47 1361 177
rect 1425 47 1455 177
rect 1509 47 1539 177
rect 1603 47 1633 177
rect 1697 47 1727 177
rect 1791 47 1821 177
<< scpmoshvt >>
rect 81 297 117 497
rect 279 297 315 497
rect 373 297 409 497
rect 467 297 503 497
rect 561 297 597 497
rect 655 297 691 497
rect 749 297 785 497
rect 843 297 879 497
rect 937 297 973 497
rect 1135 297 1171 497
rect 1229 297 1265 497
rect 1323 297 1359 497
rect 1417 297 1453 497
rect 1511 297 1547 497
rect 1605 297 1641 497
rect 1699 297 1735 497
rect 1793 297 1829 497
<< ndiff >>
rect 27 161 89 177
rect 27 127 35 161
rect 69 127 89 161
rect 27 93 89 127
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 93 171 177
rect 119 59 129 93
rect 163 59 171 93
rect 119 47 171 59
rect 225 161 287 177
rect 225 127 233 161
rect 267 127 287 161
rect 225 93 287 127
rect 225 59 233 93
rect 267 59 287 93
rect 225 47 287 59
rect 317 161 381 177
rect 317 127 327 161
rect 361 127 381 161
rect 317 47 381 127
rect 411 93 475 177
rect 411 59 421 93
rect 455 59 475 93
rect 411 47 475 59
rect 505 161 569 177
rect 505 127 515 161
rect 549 127 569 161
rect 505 47 569 127
rect 599 93 663 177
rect 599 59 609 93
rect 643 59 663 93
rect 599 47 663 59
rect 693 161 757 177
rect 693 127 703 161
rect 737 127 757 161
rect 693 47 757 127
rect 787 93 851 177
rect 787 59 797 93
rect 831 59 851 93
rect 787 47 851 59
rect 881 161 945 177
rect 881 127 891 161
rect 925 127 945 161
rect 881 47 945 127
rect 975 93 1027 177
rect 975 59 985 93
rect 1019 59 1027 93
rect 975 47 1027 59
rect 1081 93 1143 177
rect 1081 59 1089 93
rect 1123 59 1143 93
rect 1081 47 1143 59
rect 1173 161 1237 177
rect 1173 127 1183 161
rect 1217 127 1237 161
rect 1173 47 1237 127
rect 1267 93 1331 177
rect 1267 59 1277 93
rect 1311 59 1331 93
rect 1267 47 1331 59
rect 1361 161 1425 177
rect 1361 127 1371 161
rect 1405 127 1425 161
rect 1361 47 1425 127
rect 1455 161 1509 177
rect 1455 127 1465 161
rect 1499 127 1509 161
rect 1455 93 1509 127
rect 1455 59 1465 93
rect 1499 59 1509 93
rect 1455 47 1509 59
rect 1539 93 1603 177
rect 1539 59 1559 93
rect 1593 59 1603 93
rect 1539 47 1603 59
rect 1633 161 1697 177
rect 1633 127 1653 161
rect 1687 127 1697 161
rect 1633 93 1697 127
rect 1633 59 1653 93
rect 1687 59 1697 93
rect 1633 47 1697 59
rect 1727 93 1791 177
rect 1727 59 1747 93
rect 1781 59 1791 93
rect 1727 47 1791 59
rect 1821 161 1883 177
rect 1821 127 1841 161
rect 1875 127 1883 161
rect 1821 93 1883 127
rect 1821 59 1841 93
rect 1875 59 1883 93
rect 1821 47 1883 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 171 497
rect 117 451 129 485
rect 163 451 171 485
rect 117 417 171 451
rect 117 383 129 417
rect 163 383 171 417
rect 117 297 171 383
rect 225 485 279 497
rect 225 451 233 485
rect 267 451 279 485
rect 225 417 279 451
rect 225 383 233 417
rect 267 383 279 417
rect 225 349 279 383
rect 225 315 233 349
rect 267 315 279 349
rect 225 297 279 315
rect 315 485 373 497
rect 315 451 327 485
rect 361 451 373 485
rect 315 417 373 451
rect 315 383 327 417
rect 361 383 373 417
rect 315 349 373 383
rect 315 315 327 349
rect 361 315 373 349
rect 315 297 373 315
rect 409 485 467 497
rect 409 451 421 485
rect 455 451 467 485
rect 409 417 467 451
rect 409 383 421 417
rect 455 383 467 417
rect 409 297 467 383
rect 503 485 561 497
rect 503 451 515 485
rect 549 451 561 485
rect 503 417 561 451
rect 503 383 515 417
rect 549 383 561 417
rect 503 349 561 383
rect 503 315 515 349
rect 549 315 561 349
rect 503 297 561 315
rect 597 485 655 497
rect 597 451 609 485
rect 643 451 655 485
rect 597 417 655 451
rect 597 383 609 417
rect 643 383 655 417
rect 597 297 655 383
rect 691 485 749 497
rect 691 451 703 485
rect 737 451 749 485
rect 691 417 749 451
rect 691 383 703 417
rect 737 383 749 417
rect 691 349 749 383
rect 691 315 703 349
rect 737 315 749 349
rect 691 297 749 315
rect 785 485 843 497
rect 785 451 797 485
rect 831 451 843 485
rect 785 417 843 451
rect 785 383 797 417
rect 831 383 843 417
rect 785 297 843 383
rect 879 485 937 497
rect 879 451 891 485
rect 925 451 937 485
rect 879 417 937 451
rect 879 383 891 417
rect 925 383 937 417
rect 879 349 937 383
rect 879 315 891 349
rect 925 315 937 349
rect 879 297 937 315
rect 973 485 1135 497
rect 973 451 1001 485
rect 1035 451 1073 485
rect 1107 451 1135 485
rect 973 417 1135 451
rect 973 383 1001 417
rect 1035 383 1073 417
rect 1107 383 1135 417
rect 973 297 1135 383
rect 1171 485 1229 497
rect 1171 451 1183 485
rect 1217 451 1229 485
rect 1171 417 1229 451
rect 1171 383 1183 417
rect 1217 383 1229 417
rect 1171 349 1229 383
rect 1171 315 1183 349
rect 1217 315 1229 349
rect 1171 297 1229 315
rect 1265 485 1323 497
rect 1265 451 1277 485
rect 1311 451 1323 485
rect 1265 417 1323 451
rect 1265 383 1277 417
rect 1311 383 1323 417
rect 1265 297 1323 383
rect 1359 485 1417 497
rect 1359 451 1371 485
rect 1405 451 1417 485
rect 1359 417 1417 451
rect 1359 383 1371 417
rect 1405 383 1417 417
rect 1359 349 1417 383
rect 1359 315 1371 349
rect 1405 315 1417 349
rect 1359 297 1417 315
rect 1453 485 1511 497
rect 1453 451 1465 485
rect 1499 451 1511 485
rect 1453 417 1511 451
rect 1453 383 1465 417
rect 1499 383 1511 417
rect 1453 297 1511 383
rect 1547 485 1605 497
rect 1547 451 1559 485
rect 1593 451 1605 485
rect 1547 417 1605 451
rect 1547 383 1559 417
rect 1593 383 1605 417
rect 1547 349 1605 383
rect 1547 315 1559 349
rect 1593 315 1605 349
rect 1547 297 1605 315
rect 1641 485 1699 497
rect 1641 451 1653 485
rect 1687 451 1699 485
rect 1641 417 1699 451
rect 1641 383 1653 417
rect 1687 383 1699 417
rect 1641 297 1699 383
rect 1735 485 1793 497
rect 1735 451 1747 485
rect 1781 451 1793 485
rect 1735 417 1793 451
rect 1735 383 1747 417
rect 1781 383 1793 417
rect 1735 349 1793 383
rect 1735 315 1747 349
rect 1781 315 1793 349
rect 1735 297 1793 315
rect 1829 485 1883 497
rect 1829 451 1841 485
rect 1875 451 1883 485
rect 1829 417 1883 451
rect 1829 383 1841 417
rect 1875 383 1883 417
rect 1829 349 1883 383
rect 1829 315 1841 349
rect 1875 315 1883 349
rect 1829 297 1883 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 59 163 93
rect 233 127 267 161
rect 233 59 267 93
rect 327 127 361 161
rect 421 59 455 93
rect 515 127 549 161
rect 609 59 643 93
rect 703 127 737 161
rect 797 59 831 93
rect 891 127 925 161
rect 985 59 1019 93
rect 1089 59 1123 93
rect 1183 127 1217 161
rect 1277 59 1311 93
rect 1371 127 1405 161
rect 1465 127 1499 161
rect 1465 59 1499 93
rect 1559 59 1593 93
rect 1653 127 1687 161
rect 1653 59 1687 93
rect 1747 59 1781 93
rect 1841 127 1875 161
rect 1841 59 1875 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 233 451 267 485
rect 233 383 267 417
rect 233 315 267 349
rect 327 451 361 485
rect 327 383 361 417
rect 327 315 361 349
rect 421 451 455 485
rect 421 383 455 417
rect 515 451 549 485
rect 515 383 549 417
rect 515 315 549 349
rect 609 451 643 485
rect 609 383 643 417
rect 703 451 737 485
rect 703 383 737 417
rect 703 315 737 349
rect 797 451 831 485
rect 797 383 831 417
rect 891 451 925 485
rect 891 383 925 417
rect 891 315 925 349
rect 1001 451 1035 485
rect 1073 451 1107 485
rect 1001 383 1035 417
rect 1073 383 1107 417
rect 1183 451 1217 485
rect 1183 383 1217 417
rect 1183 315 1217 349
rect 1277 451 1311 485
rect 1277 383 1311 417
rect 1371 451 1405 485
rect 1371 383 1405 417
rect 1371 315 1405 349
rect 1465 451 1499 485
rect 1465 383 1499 417
rect 1559 451 1593 485
rect 1559 383 1593 417
rect 1559 315 1593 349
rect 1653 451 1687 485
rect 1653 383 1687 417
rect 1747 451 1781 485
rect 1747 383 1781 417
rect 1747 315 1781 349
rect 1841 451 1875 485
rect 1841 383 1875 417
rect 1841 315 1875 349
<< poly >>
rect 81 497 117 523
rect 279 497 315 523
rect 373 497 409 523
rect 467 497 503 523
rect 561 497 597 523
rect 655 497 691 523
rect 749 497 785 523
rect 843 497 879 523
rect 937 497 973 523
rect 1135 497 1171 523
rect 1229 497 1265 523
rect 1323 497 1359 523
rect 1417 497 1453 523
rect 1511 497 1547 523
rect 1605 497 1641 523
rect 1699 497 1735 523
rect 1793 497 1829 523
rect 81 282 117 297
rect 279 282 315 297
rect 373 282 409 297
rect 467 282 503 297
rect 561 282 597 297
rect 655 282 691 297
rect 749 282 785 297
rect 843 282 879 297
rect 937 282 973 297
rect 1135 282 1171 297
rect 1229 282 1265 297
rect 1323 282 1359 297
rect 1417 282 1453 297
rect 1511 282 1547 297
rect 1605 282 1641 297
rect 1699 282 1735 297
rect 1793 282 1829 297
rect 79 265 119 282
rect 76 261 119 265
rect 22 249 119 261
rect 277 259 317 282
rect 371 259 411 282
rect 465 259 505 282
rect 559 259 599 282
rect 653 259 693 282
rect 747 259 787 282
rect 841 259 881 282
rect 935 261 975 282
rect 935 259 1008 261
rect 1133 259 1173 282
rect 1227 259 1267 282
rect 1321 259 1361 282
rect 1415 259 1455 282
rect 22 215 38 249
rect 72 215 119 249
rect 22 203 119 215
rect 211 249 599 259
rect 211 215 227 249
rect 261 215 327 249
rect 361 215 599 249
rect 211 205 599 215
rect 641 249 1008 259
rect 641 215 657 249
rect 691 215 763 249
rect 797 215 858 249
rect 892 215 948 249
rect 982 215 1008 249
rect 641 205 1008 215
rect 1054 249 1455 259
rect 1054 215 1070 249
rect 1104 215 1183 249
rect 1217 215 1277 249
rect 1311 215 1372 249
rect 1406 215 1455 249
rect 1054 205 1455 215
rect 89 177 119 203
rect 287 177 317 205
rect 381 177 411 205
rect 475 177 505 205
rect 569 177 599 205
rect 663 177 693 205
rect 757 177 787 205
rect 851 177 881 205
rect 945 203 1008 205
rect 945 177 975 203
rect 1143 177 1173 205
rect 1237 177 1267 205
rect 1331 177 1361 205
rect 1425 177 1455 205
rect 1509 259 1549 282
rect 1603 259 1643 282
rect 1697 259 1737 282
rect 1791 261 1831 282
rect 1791 259 1897 261
rect 1509 249 1897 259
rect 1509 215 1559 249
rect 1593 215 1653 249
rect 1687 215 1747 249
rect 1781 215 1847 249
rect 1881 215 1897 249
rect 1509 205 1897 215
rect 1509 177 1539 205
rect 1603 177 1633 205
rect 1697 177 1727 205
rect 1791 203 1897 205
rect 1791 177 1821 203
rect 89 21 119 47
rect 287 21 317 47
rect 381 21 411 47
rect 475 21 505 47
rect 569 21 599 47
rect 663 21 693 47
rect 757 21 787 47
rect 851 21 881 47
rect 945 21 975 47
rect 1143 21 1173 47
rect 1237 21 1267 47
rect 1331 21 1361 47
rect 1425 21 1455 47
rect 1509 21 1539 47
rect 1603 21 1633 47
rect 1697 21 1727 47
rect 1791 21 1821 47
<< polycont >>
rect 38 215 72 249
rect 227 215 261 249
rect 327 215 361 249
rect 657 215 691 249
rect 763 215 797 249
rect 858 215 892 249
rect 948 215 982 249
rect 1070 215 1104 249
rect 1183 215 1217 249
rect 1277 215 1311 249
rect 1372 215 1406 249
rect 1559 215 1593 249
rect 1653 215 1687 249
rect 1747 215 1781 249
rect 1847 215 1881 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 18 485 85 493
rect 18 451 35 485
rect 69 451 85 485
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 18 349 85 383
rect 129 485 267 527
rect 163 451 233 485
rect 129 417 267 451
rect 163 383 233 417
rect 129 367 267 383
rect 18 315 35 349
rect 69 333 85 349
rect 209 349 267 367
rect 69 315 171 333
rect 18 299 171 315
rect 209 315 233 349
rect 209 299 267 315
rect 301 485 377 493
rect 301 451 327 485
rect 361 451 377 485
rect 301 417 377 451
rect 301 383 327 417
rect 361 383 377 417
rect 301 349 377 383
rect 421 485 455 527
rect 421 417 455 451
rect 421 367 455 383
rect 489 485 565 493
rect 489 451 515 485
rect 549 451 565 485
rect 489 417 565 451
rect 489 383 515 417
rect 549 383 565 417
rect 301 315 327 349
rect 361 333 377 349
rect 489 349 565 383
rect 609 485 643 527
rect 609 417 643 451
rect 609 367 643 383
rect 677 485 753 493
rect 677 451 703 485
rect 737 451 753 485
rect 677 417 753 451
rect 677 383 703 417
rect 737 383 753 417
rect 489 333 515 349
rect 361 315 515 333
rect 549 333 565 349
rect 677 349 753 383
rect 797 485 831 527
rect 797 417 831 451
rect 797 367 831 383
rect 865 485 941 493
rect 865 451 891 485
rect 925 451 941 485
rect 865 417 941 451
rect 865 383 891 417
rect 925 383 941 417
rect 677 333 703 349
rect 549 315 703 333
rect 737 333 753 349
rect 865 349 941 383
rect 985 485 1123 527
rect 985 451 1001 485
rect 1035 451 1073 485
rect 1107 451 1123 485
rect 985 417 1123 451
rect 985 383 1001 417
rect 1035 383 1073 417
rect 1107 383 1123 417
rect 985 367 1123 383
rect 1157 485 1233 493
rect 1157 451 1183 485
rect 1217 451 1233 485
rect 1157 417 1233 451
rect 1157 383 1183 417
rect 1217 383 1233 417
rect 865 333 891 349
rect 737 315 891 333
rect 925 333 941 349
rect 1157 349 1233 383
rect 1277 485 1311 527
rect 1277 417 1311 451
rect 1277 367 1311 383
rect 1345 485 1421 493
rect 1345 451 1371 485
rect 1405 451 1421 485
rect 1345 417 1421 451
rect 1345 383 1371 417
rect 1405 383 1421 417
rect 1157 333 1183 349
rect 925 315 1183 333
rect 1217 333 1233 349
rect 1345 349 1421 383
rect 1465 485 1499 527
rect 1465 417 1499 451
rect 1465 367 1499 383
rect 1533 485 1609 493
rect 1533 451 1559 485
rect 1593 451 1609 485
rect 1533 417 1609 451
rect 1533 383 1559 417
rect 1593 383 1609 417
rect 1345 333 1371 349
rect 1217 315 1371 333
rect 1405 333 1421 349
rect 1533 349 1609 383
rect 1653 485 1687 527
rect 1653 417 1687 451
rect 1653 367 1687 383
rect 1721 485 1797 493
rect 1721 451 1747 485
rect 1781 451 1797 485
rect 1721 417 1797 451
rect 1721 383 1747 417
rect 1781 383 1797 417
rect 1533 333 1559 349
rect 1405 315 1559 333
rect 1593 333 1609 349
rect 1721 349 1797 383
rect 1721 333 1747 349
rect 1593 315 1747 333
rect 1781 315 1797 349
rect 132 255 171 299
rect 301 289 1797 315
rect 1841 485 1892 527
rect 1875 451 1892 485
rect 1841 417 1892 451
rect 1875 383 1892 417
rect 1841 349 1892 383
rect 1875 315 1892 349
rect 1841 289 1892 315
rect 22 249 88 255
rect 22 215 38 249
rect 72 215 88 249
rect 132 249 395 255
rect 132 215 227 249
rect 261 215 327 249
rect 361 215 395 249
rect 132 181 171 215
rect 482 181 568 289
rect 636 249 1008 255
rect 636 215 657 249
rect 691 215 763 249
rect 797 215 858 249
rect 892 215 948 249
rect 982 215 1008 249
rect 1048 249 1422 255
rect 1048 215 1070 249
rect 1104 215 1183 249
rect 1217 215 1277 249
rect 1311 215 1372 249
rect 1406 215 1422 249
rect 1533 249 1901 255
rect 1533 215 1559 249
rect 1593 215 1653 249
rect 1687 215 1747 249
rect 1781 215 1847 249
rect 1881 215 1901 249
rect 18 161 171 181
rect 18 127 35 161
rect 69 147 171 161
rect 217 161 267 181
rect 69 127 85 147
rect 18 93 85 127
rect 217 127 233 161
rect 301 161 568 181
rect 301 127 327 161
rect 361 127 515 161
rect 549 127 568 161
rect 677 161 1421 181
rect 677 127 703 161
rect 737 127 891 161
rect 925 127 1183 161
rect 1217 127 1371 161
rect 1405 127 1421 161
rect 1465 161 1892 181
rect 1499 147 1653 161
rect 1499 127 1515 147
rect 18 59 35 93
rect 69 59 85 93
rect 18 51 85 59
rect 129 93 179 109
rect 163 59 179 93
rect 129 17 179 59
rect 217 93 267 127
rect 1465 93 1515 127
rect 1627 127 1653 147
rect 1687 147 1841 161
rect 1687 127 1703 147
rect 217 59 233 93
rect 267 59 421 93
rect 455 59 609 93
rect 643 59 797 93
rect 831 59 985 93
rect 1019 59 1035 93
rect 217 51 1035 59
rect 1073 59 1089 93
rect 1123 59 1277 93
rect 1311 59 1465 93
rect 1499 59 1515 93
rect 1073 51 1515 59
rect 1559 93 1593 109
rect 1559 17 1593 59
rect 1627 93 1703 127
rect 1815 127 1841 147
rect 1875 127 1892 161
rect 1627 59 1653 93
rect 1687 59 1703 93
rect 1627 51 1703 59
rect 1747 93 1781 109
rect 1747 17 1781 59
rect 1815 93 1892 127
rect 1815 59 1841 93
rect 1875 59 1892 93
rect 1815 51 1892 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 1325 221 1369 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 1683 221 1717 255 0 FreeSans 250 0 0 0 D
port 4 nsew signal input
flabel locali s 1594 221 1628 255 0 FreeSans 250 0 0 0 D
port 4 nsew signal input
flabel locali s 1762 221 1796 255 0 FreeSans 250 0 0 0 D
port 4 nsew signal input
flabel locali s 1140 221 1184 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 1048 221 1082 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 948 221 982 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 858 221 892 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 764 221 798 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 677 221 711 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 534 153 568 187 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 534 221 568 255 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 534 289 568 323 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel locali s 1242 221 1286 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 1855 221 1889 255 0 FreeSans 250 0 0 0 D
port 4 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_END 1636080
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1620730
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
