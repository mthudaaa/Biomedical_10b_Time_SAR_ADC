magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 335 157 1287 203
rect 1 21 1287 157
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 131
rect 183 47 213 131
rect 423 47 453 177
rect 517 47 547 177
rect 611 47 641 177
rect 705 47 735 177
rect 897 47 927 177
rect 991 47 1021 177
rect 1085 47 1115 177
rect 1179 47 1209 177
<< scpmoshvt >>
rect 81 413 117 497
rect 175 413 211 497
rect 415 297 451 497
rect 509 297 545 497
rect 603 297 639 497
rect 697 297 733 497
rect 889 297 925 497
rect 983 297 1019 497
rect 1077 297 1113 497
rect 1171 297 1207 497
<< ndiff >>
rect 27 109 89 131
rect 27 75 35 109
rect 69 75 89 109
rect 27 47 89 75
rect 119 93 183 131
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 109 307 131
rect 213 75 223 109
rect 257 75 307 109
rect 213 47 307 75
rect 361 101 423 177
rect 361 67 369 101
rect 403 67 423 101
rect 361 47 423 67
rect 453 165 517 177
rect 453 131 463 165
rect 497 131 517 165
rect 453 47 517 131
rect 547 97 611 177
rect 547 63 557 97
rect 591 63 611 97
rect 547 47 611 63
rect 641 165 705 177
rect 641 131 651 165
rect 685 131 705 165
rect 641 47 705 131
rect 735 97 787 177
rect 735 63 745 97
rect 779 63 787 97
rect 735 47 787 63
rect 841 97 897 177
rect 841 63 849 97
rect 883 63 897 97
rect 841 47 897 63
rect 927 165 991 177
rect 927 131 937 165
rect 971 131 991 165
rect 927 47 991 131
rect 1021 165 1085 177
rect 1021 131 1031 165
rect 1065 131 1085 165
rect 1021 97 1085 131
rect 1021 63 1031 97
rect 1065 63 1085 97
rect 1021 47 1085 63
rect 1115 97 1179 177
rect 1115 63 1125 97
rect 1159 63 1179 97
rect 1115 47 1179 63
rect 1209 165 1261 177
rect 1209 131 1219 165
rect 1253 131 1261 165
rect 1209 97 1261 131
rect 1209 63 1219 97
rect 1253 63 1261 97
rect 1209 47 1261 63
<< pdiff >>
rect 27 472 81 497
rect 27 438 35 472
rect 69 438 81 472
rect 27 413 81 438
rect 117 489 175 497
rect 117 455 129 489
rect 163 455 175 489
rect 117 413 175 455
rect 211 483 307 497
rect 211 449 223 483
rect 257 449 307 483
rect 211 413 307 449
rect 361 485 415 497
rect 361 451 369 485
rect 403 451 415 485
rect 361 417 415 451
rect 361 383 369 417
rect 403 383 415 417
rect 361 349 415 383
rect 361 315 369 349
rect 403 315 415 349
rect 361 297 415 315
rect 451 477 509 497
rect 451 443 463 477
rect 497 443 509 477
rect 451 374 509 443
rect 451 340 463 374
rect 497 340 509 374
rect 451 297 509 340
rect 545 485 603 497
rect 545 451 557 485
rect 591 451 603 485
rect 545 417 603 451
rect 545 383 557 417
rect 591 383 603 417
rect 545 297 603 383
rect 639 485 697 497
rect 639 451 651 485
rect 685 451 697 485
rect 639 417 697 451
rect 639 383 651 417
rect 685 383 697 417
rect 639 349 697 383
rect 639 315 651 349
rect 685 315 697 349
rect 639 297 697 315
rect 733 485 889 497
rect 733 451 761 485
rect 795 451 833 485
rect 867 451 889 485
rect 733 417 889 451
rect 733 383 761 417
rect 795 383 833 417
rect 867 383 889 417
rect 733 297 889 383
rect 925 485 983 497
rect 925 451 937 485
rect 971 451 983 485
rect 925 417 983 451
rect 925 383 937 417
rect 971 383 983 417
rect 925 349 983 383
rect 925 315 937 349
rect 971 315 983 349
rect 925 297 983 315
rect 1019 485 1077 497
rect 1019 451 1031 485
rect 1065 451 1077 485
rect 1019 417 1077 451
rect 1019 383 1031 417
rect 1065 383 1077 417
rect 1019 297 1077 383
rect 1113 485 1171 497
rect 1113 451 1125 485
rect 1159 451 1171 485
rect 1113 417 1171 451
rect 1113 383 1125 417
rect 1159 383 1171 417
rect 1113 349 1171 383
rect 1113 315 1125 349
rect 1159 315 1171 349
rect 1113 297 1171 315
rect 1207 485 1261 497
rect 1207 451 1219 485
rect 1253 451 1261 485
rect 1207 417 1261 451
rect 1207 383 1219 417
rect 1253 383 1261 417
rect 1207 349 1261 383
rect 1207 315 1219 349
rect 1253 315 1261 349
rect 1207 297 1261 315
<< ndiffc >>
rect 35 75 69 109
rect 129 59 163 93
rect 223 75 257 109
rect 369 67 403 101
rect 463 131 497 165
rect 557 63 591 97
rect 651 131 685 165
rect 745 63 779 97
rect 849 63 883 97
rect 937 131 971 165
rect 1031 131 1065 165
rect 1031 63 1065 97
rect 1125 63 1159 97
rect 1219 131 1253 165
rect 1219 63 1253 97
<< pdiffc >>
rect 35 438 69 472
rect 129 455 163 489
rect 223 449 257 483
rect 369 451 403 485
rect 369 383 403 417
rect 369 315 403 349
rect 463 443 497 477
rect 463 340 497 374
rect 557 451 591 485
rect 557 383 591 417
rect 651 451 685 485
rect 651 383 685 417
rect 651 315 685 349
rect 761 451 795 485
rect 833 451 867 485
rect 761 383 795 417
rect 833 383 867 417
rect 937 451 971 485
rect 937 383 971 417
rect 937 315 971 349
rect 1031 451 1065 485
rect 1031 383 1065 417
rect 1125 451 1159 485
rect 1125 383 1159 417
rect 1125 315 1159 349
rect 1219 451 1253 485
rect 1219 383 1253 417
rect 1219 315 1253 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 415 497 451 523
rect 509 497 545 523
rect 603 497 639 523
rect 697 497 733 523
rect 889 497 925 523
rect 983 497 1019 523
rect 1077 497 1113 523
rect 1171 497 1207 523
rect 81 398 117 413
rect 175 398 211 413
rect 79 387 119 398
rect 46 357 119 387
rect 46 280 76 357
rect 173 284 213 398
rect 21 264 76 280
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 128 268 213 284
rect 415 282 451 297
rect 509 282 545 297
rect 603 282 639 297
rect 697 282 733 297
rect 889 282 925 297
rect 983 282 1019 297
rect 1077 282 1113 297
rect 1171 282 1207 297
rect 128 234 138 268
rect 172 234 213 268
rect 413 265 453 282
rect 128 218 213 234
rect 46 176 76 214
rect 46 146 119 176
rect 89 131 119 146
rect 183 131 213 218
rect 290 259 453 265
rect 507 259 547 282
rect 601 259 641 282
rect 695 259 735 282
rect 290 249 547 259
rect 290 215 300 249
rect 334 215 547 249
rect 290 205 547 215
rect 589 249 735 259
rect 589 215 605 249
rect 639 215 735 249
rect 589 205 735 215
rect 290 199 453 205
rect 423 177 453 199
rect 517 177 547 205
rect 611 177 641 205
rect 705 177 735 205
rect 887 259 927 282
rect 981 259 1021 282
rect 1075 259 1115 282
rect 1169 261 1209 282
rect 1169 259 1248 261
rect 887 249 1021 259
rect 887 215 937 249
rect 971 215 1021 249
rect 887 205 1021 215
rect 1063 249 1248 259
rect 1063 215 1079 249
rect 1113 215 1198 249
rect 1232 215 1248 249
rect 1063 205 1248 215
rect 887 203 927 205
rect 897 177 927 203
rect 991 177 1021 205
rect 1085 177 1115 205
rect 1179 203 1248 205
rect 1179 177 1209 203
rect 89 21 119 47
rect 183 21 213 47
rect 423 21 453 47
rect 517 21 547 47
rect 611 21 641 47
rect 705 21 735 47
rect 897 21 927 47
rect 991 21 1021 47
rect 1085 21 1115 47
rect 1179 21 1209 47
<< polycont >>
rect 32 230 66 264
rect 138 234 172 268
rect 300 215 334 249
rect 605 215 639 249
rect 937 215 971 249
rect 1079 215 1113 249
rect 1198 215 1232 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 108 489 163 527
rect 17 472 74 488
rect 17 438 35 472
rect 69 438 74 472
rect 108 455 129 489
rect 108 439 163 455
rect 197 483 335 493
rect 197 449 223 483
rect 257 449 335 483
rect 17 396 74 438
rect 197 430 335 449
rect 17 357 266 396
rect 17 264 66 323
rect 17 230 32 264
rect 17 214 66 230
rect 112 268 188 323
rect 112 234 138 268
rect 172 234 188 268
rect 112 214 188 234
rect 232 255 266 357
rect 232 180 266 221
rect 17 146 266 180
rect 300 249 335 430
rect 369 485 403 527
rect 369 417 403 451
rect 369 349 403 383
rect 369 299 403 315
rect 437 477 497 493
rect 437 443 463 477
rect 437 374 497 443
rect 437 340 463 374
rect 531 485 591 527
rect 531 451 557 485
rect 531 417 591 451
rect 531 383 557 417
rect 531 367 591 383
rect 625 485 701 493
rect 625 451 651 485
rect 685 451 701 485
rect 625 417 701 451
rect 625 383 651 417
rect 685 383 701 417
rect 437 333 497 340
rect 625 349 701 383
rect 745 485 877 527
rect 745 451 761 485
rect 795 451 833 485
rect 867 451 877 485
rect 745 417 877 451
rect 745 383 761 417
rect 795 383 833 417
rect 867 383 877 417
rect 745 367 877 383
rect 911 485 987 493
rect 911 451 937 485
rect 971 451 987 485
rect 911 417 987 451
rect 911 383 937 417
rect 971 383 987 417
rect 625 333 651 349
rect 437 315 651 333
rect 685 333 701 349
rect 911 349 987 383
rect 1031 485 1065 527
rect 1031 417 1065 451
rect 1031 367 1065 383
rect 1099 485 1175 493
rect 1099 451 1125 485
rect 1159 451 1175 485
rect 1099 417 1175 451
rect 1099 383 1125 417
rect 1159 383 1175 417
rect 911 333 937 349
rect 685 315 937 333
rect 971 333 987 349
rect 1099 349 1175 383
rect 1099 333 1125 349
rect 971 315 1125 333
rect 1159 315 1175 349
rect 334 215 335 249
rect 17 109 69 146
rect 300 112 335 215
rect 437 289 1175 315
rect 1219 485 1269 527
rect 1253 451 1269 485
rect 1219 417 1269 451
rect 1253 383 1269 417
rect 1219 349 1269 383
rect 1253 315 1269 349
rect 1219 289 1269 315
rect 437 165 526 289
rect 589 249 631 255
rect 589 215 605 249
rect 639 215 665 221
rect 699 215 809 289
rect 848 249 990 255
rect 848 215 937 249
rect 971 215 990 249
rect 1063 249 1259 255
rect 1063 215 1079 249
rect 1113 215 1198 249
rect 1232 215 1259 249
rect 437 131 463 165
rect 497 131 526 165
rect 625 165 987 181
rect 625 131 651 165
rect 685 131 937 165
rect 971 131 987 165
rect 1031 165 1269 181
rect 1065 147 1219 165
rect 1065 131 1081 147
rect 197 109 335 112
rect 17 75 35 109
rect 17 51 69 75
rect 103 93 163 109
rect 103 59 129 93
rect 103 17 163 59
rect 197 75 223 109
rect 257 75 335 109
rect 197 51 335 75
rect 369 101 403 117
rect 1031 97 1081 131
rect 1193 131 1219 147
rect 1253 131 1269 165
rect 403 67 557 97
rect 369 63 557 67
rect 591 63 745 97
rect 779 63 795 97
rect 369 51 795 63
rect 833 63 849 97
rect 883 63 1031 97
rect 1065 63 1081 97
rect 833 51 1081 63
rect 1125 97 1159 113
rect 1125 17 1159 63
rect 1193 97 1269 131
rect 1193 63 1219 97
rect 1253 63 1269 97
rect 1193 51 1269 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 232 221 266 255
rect 631 249 665 255
rect 631 221 639 249
rect 639 221 665 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 220 255 677 261
rect 220 221 232 255
rect 266 221 631 255
rect 665 221 677 255
rect 220 215 677 221
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 1129 221 1163 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 1210 221 1244 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 948 221 982 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel locali s 132 289 166 323 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 132 221 166 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 762 289 796 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 758 221 792 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 858 221 892 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4bb_2
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 1654128
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1643532
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
