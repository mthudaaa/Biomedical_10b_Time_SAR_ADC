magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 1255 157 1444 201
rect 1790 157 2080 203
rect 1 145 895 157
rect 1113 145 2080 157
rect 1 21 2080 145
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 173 47 203 131
rect 387 47 417 131
rect 477 47 507 131
rect 585 47 615 131
rect 691 47 721 131
rect 767 47 797 131
rect 981 47 1011 119
rect 1087 47 1117 119
rect 1189 47 1219 131
rect 1338 47 1368 175
rect 1446 47 1476 119
rect 1551 47 1581 119
rect 1647 47 1677 131
rect 1878 47 1908 177
rect 1962 47 1992 177
<< scpmoshvt >>
rect 82 363 118 491
rect 176 363 212 491
rect 374 369 410 497
rect 468 369 504 497
rect 572 369 608 497
rect 666 369 702 497
rect 769 369 805 497
rect 982 413 1018 497
rect 1085 413 1121 497
rect 1191 413 1227 497
rect 1330 347 1366 497
rect 1438 413 1474 497
rect 1534 413 1570 497
rect 1649 413 1685 497
rect 1870 297 1906 497
rect 1964 297 2000 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 173 131
rect 109 59 129 93
rect 163 59 173 93
rect 109 47 173 59
rect 203 119 265 131
rect 203 85 223 119
rect 257 85 265 119
rect 203 47 265 85
rect 319 89 387 131
rect 319 55 331 89
rect 365 55 387 89
rect 319 47 387 55
rect 417 89 477 131
rect 417 55 431 89
rect 465 55 477 89
rect 417 47 477 55
rect 507 47 585 131
rect 615 89 691 131
rect 615 55 636 89
rect 670 55 691 89
rect 615 47 691 55
rect 721 47 767 131
rect 797 89 869 131
rect 1281 131 1338 175
rect 1139 119 1189 131
rect 797 55 823 89
rect 857 55 869 89
rect 797 47 869 55
rect 925 107 981 119
rect 925 73 933 107
rect 967 73 981 107
rect 925 47 981 73
rect 1011 107 1087 119
rect 1011 73 1043 107
rect 1077 73 1087 107
rect 1011 47 1087 73
rect 1117 47 1189 119
rect 1219 101 1338 131
rect 1219 67 1279 101
rect 1313 67 1338 101
rect 1219 47 1338 67
rect 1368 119 1418 175
rect 1816 162 1878 177
rect 1597 119 1647 131
rect 1368 107 1446 119
rect 1368 73 1402 107
rect 1436 73 1446 107
rect 1368 47 1446 73
rect 1476 107 1551 119
rect 1476 73 1507 107
rect 1541 73 1551 107
rect 1476 47 1551 73
rect 1581 47 1647 119
rect 1677 107 1762 131
rect 1677 73 1720 107
rect 1754 73 1762 107
rect 1677 47 1762 73
rect 1816 128 1824 162
rect 1858 128 1878 162
rect 1816 94 1878 128
rect 1816 60 1824 94
rect 1858 60 1878 94
rect 1816 47 1878 60
rect 1908 123 1962 177
rect 1908 89 1918 123
rect 1952 89 1962 123
rect 1908 47 1962 89
rect 1992 164 2054 177
rect 1992 130 2012 164
rect 2046 130 2054 164
rect 1992 96 2054 130
rect 1992 62 2012 96
rect 2046 62 2054 96
rect 1992 47 2054 62
<< pdiff >>
rect 28 477 82 491
rect 28 443 36 477
rect 70 443 82 477
rect 28 409 82 443
rect 28 375 36 409
rect 70 375 82 409
rect 28 363 82 375
rect 118 461 176 491
rect 118 427 130 461
rect 164 427 176 461
rect 118 363 176 427
rect 212 477 266 491
rect 212 443 224 477
rect 258 443 266 477
rect 212 409 266 443
rect 212 375 224 409
rect 258 375 266 409
rect 212 363 266 375
rect 320 452 374 497
rect 320 418 328 452
rect 362 418 374 452
rect 320 369 374 418
rect 410 483 468 497
rect 410 449 422 483
rect 456 449 468 483
rect 410 369 468 449
rect 504 369 572 497
rect 608 483 666 497
rect 608 449 620 483
rect 654 449 666 483
rect 608 369 666 449
rect 702 369 769 497
rect 805 483 864 497
rect 805 449 822 483
rect 856 449 864 483
rect 805 369 864 449
rect 918 472 982 497
rect 918 438 926 472
rect 960 438 982 472
rect 918 413 982 438
rect 1018 472 1085 497
rect 1018 438 1035 472
rect 1069 438 1085 472
rect 1018 413 1085 438
rect 1121 413 1191 497
rect 1227 485 1330 497
rect 1227 451 1280 485
rect 1314 451 1330 485
rect 1227 417 1330 451
rect 1227 413 1280 417
rect 1244 383 1280 413
rect 1314 383 1330 417
rect 1244 347 1330 383
rect 1366 477 1438 497
rect 1366 443 1378 477
rect 1412 443 1438 477
rect 1366 413 1438 443
rect 1474 467 1534 497
rect 1474 433 1486 467
rect 1520 433 1534 467
rect 1474 413 1534 433
rect 1570 413 1649 497
rect 1685 477 1762 497
rect 1685 443 1719 477
rect 1753 443 1762 477
rect 1685 413 1762 443
rect 1816 475 1870 497
rect 1816 441 1824 475
rect 1858 441 1870 475
rect 1366 347 1421 413
rect 1816 407 1870 441
rect 1816 373 1824 407
rect 1858 373 1870 407
rect 1816 297 1870 373
rect 1906 455 1964 497
rect 1906 421 1918 455
rect 1952 421 1964 455
rect 1906 375 1964 421
rect 1906 341 1918 375
rect 1952 341 1964 375
rect 1906 297 1964 341
rect 2000 479 2054 497
rect 2000 445 2012 479
rect 2046 445 2054 479
rect 2000 411 2054 445
rect 2000 377 2012 411
rect 2046 377 2054 411
rect 2000 343 2054 377
rect 2000 309 2012 343
rect 2046 309 2054 343
rect 2000 297 2054 309
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 331 55 365 89
rect 431 55 465 89
rect 636 55 670 89
rect 823 55 857 89
rect 933 73 967 107
rect 1043 73 1077 107
rect 1279 67 1313 101
rect 1402 73 1436 107
rect 1507 73 1541 107
rect 1720 73 1754 107
rect 1824 128 1858 162
rect 1824 60 1858 94
rect 1918 89 1952 123
rect 2012 130 2046 164
rect 2012 62 2046 96
<< pdiffc >>
rect 36 443 70 477
rect 36 375 70 409
rect 130 427 164 461
rect 224 443 258 477
rect 224 375 258 409
rect 328 418 362 452
rect 422 449 456 483
rect 620 449 654 483
rect 822 449 856 483
rect 926 438 960 472
rect 1035 438 1069 472
rect 1280 451 1314 485
rect 1280 383 1314 417
rect 1378 443 1412 477
rect 1486 433 1520 467
rect 1719 443 1753 477
rect 1824 441 1858 475
rect 1824 373 1858 407
rect 1918 421 1952 455
rect 1918 341 1952 375
rect 2012 445 2046 479
rect 2012 377 2046 411
rect 2012 309 2046 343
<< poly >>
rect 82 491 118 517
rect 176 491 212 517
rect 374 497 410 523
rect 468 497 504 523
rect 572 497 608 523
rect 666 497 702 523
rect 769 497 805 523
rect 982 497 1018 523
rect 1085 497 1121 523
rect 1191 497 1227 523
rect 1330 497 1366 523
rect 1438 497 1474 523
rect 1534 497 1570 523
rect 1649 497 1685 523
rect 1870 497 1906 523
rect 1964 497 2000 523
rect 982 398 1018 413
rect 1085 398 1121 413
rect 1191 398 1227 413
rect 980 375 1020 398
rect 1083 381 1123 398
rect 82 348 118 363
rect 176 348 212 363
rect 374 354 410 369
rect 468 354 504 369
rect 572 354 608 369
rect 666 354 702 369
rect 769 354 805 369
rect 965 365 1041 375
rect 47 318 120 348
rect 47 265 77 318
rect 174 274 214 348
rect 372 331 412 354
rect 466 331 506 354
rect 570 337 610 354
rect 664 337 704 354
rect 372 321 506 331
rect 372 287 388 321
rect 422 301 506 321
rect 549 321 615 337
rect 422 287 438 301
rect 372 277 438 287
rect 549 287 565 321
rect 599 287 615 321
rect 549 277 615 287
rect 23 249 77 265
rect 23 215 33 249
rect 67 215 77 249
rect 129 264 214 274
rect 129 230 145 264
rect 179 230 214 264
rect 129 220 214 230
rect 23 199 77 215
rect 47 176 77 199
rect 47 146 109 176
rect 79 131 109 146
rect 173 131 203 220
rect 387 131 417 277
rect 477 225 543 235
rect 477 191 493 225
rect 527 191 543 225
rect 477 175 543 191
rect 477 131 507 175
rect 585 131 615 277
rect 664 321 718 337
rect 664 287 674 321
rect 708 287 718 321
rect 664 271 718 287
rect 767 304 807 354
rect 965 331 981 365
rect 1015 331 1041 365
rect 965 321 1041 331
rect 1083 365 1147 381
rect 1083 331 1093 365
rect 1127 331 1147 365
rect 1083 315 1147 331
rect 767 288 831 304
rect 767 254 777 288
rect 811 254 831 288
rect 1083 279 1123 315
rect 767 238 831 254
rect 981 249 1123 279
rect 657 207 721 223
rect 657 173 667 207
rect 701 173 721 207
rect 657 157 721 173
rect 691 131 721 157
rect 767 131 797 238
rect 981 119 1011 249
rect 1189 213 1229 398
rect 1438 398 1474 413
rect 1534 398 1570 413
rect 1649 398 1685 413
rect 1330 332 1366 347
rect 1328 309 1368 332
rect 1271 299 1368 309
rect 1271 265 1287 299
rect 1321 265 1368 299
rect 1271 255 1368 265
rect 1063 191 1117 207
rect 1063 157 1073 191
rect 1107 157 1117 191
rect 1063 141 1117 157
rect 1087 119 1117 141
rect 1189 203 1259 213
rect 1189 169 1209 203
rect 1243 169 1259 203
rect 1338 175 1368 255
rect 1436 315 1476 398
rect 1532 375 1572 398
rect 1647 381 1687 398
rect 1532 365 1598 375
rect 1532 331 1548 365
rect 1582 331 1598 365
rect 1532 321 1598 331
rect 1647 365 1735 381
rect 1647 331 1691 365
rect 1725 331 1735 365
rect 1647 315 1735 331
rect 1436 299 1490 315
rect 1436 265 1446 299
rect 1480 279 1490 299
rect 1480 265 1581 279
rect 1436 249 1581 265
rect 1446 191 1500 207
rect 1189 159 1259 169
rect 1189 131 1219 159
rect 1446 157 1456 191
rect 1490 157 1500 191
rect 1446 141 1500 157
rect 1446 119 1476 141
rect 1551 119 1581 249
rect 1647 131 1677 315
rect 1870 282 1906 297
rect 1964 282 2000 297
rect 1868 265 1908 282
rect 1766 249 1908 265
rect 1766 215 1776 249
rect 1810 215 1908 249
rect 1766 199 1908 215
rect 1878 177 1908 199
rect 1962 265 2002 282
rect 1962 249 2016 265
rect 1962 215 1972 249
rect 2006 215 2016 249
rect 1962 199 2016 215
rect 1962 177 1992 199
rect 79 21 109 47
rect 173 21 203 47
rect 387 21 417 47
rect 477 21 507 47
rect 585 21 615 47
rect 691 21 721 47
rect 767 21 797 47
rect 981 21 1011 47
rect 1087 21 1117 47
rect 1189 21 1219 47
rect 1338 21 1368 47
rect 1446 21 1476 47
rect 1551 21 1581 47
rect 1647 21 1677 47
rect 1878 21 1908 47
rect 1962 21 1992 47
<< polycont >>
rect 388 287 422 321
rect 565 287 599 321
rect 33 215 67 249
rect 145 230 179 264
rect 493 191 527 225
rect 674 287 708 321
rect 981 331 1015 365
rect 1093 331 1127 365
rect 777 254 811 288
rect 667 173 701 207
rect 1287 265 1321 299
rect 1073 157 1107 191
rect 1209 169 1243 203
rect 1548 331 1582 365
rect 1691 331 1725 365
rect 1446 265 1480 299
rect 1456 157 1490 191
rect 1776 215 1810 249
rect 1972 215 2006 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 36 477 70 493
rect 36 409 70 443
rect 104 461 180 527
rect 104 427 130 461
rect 164 427 180 461
rect 223 477 269 493
rect 223 443 224 477
rect 258 443 269 477
rect 223 409 269 443
rect 70 382 179 393
rect 70 375 133 382
rect 36 359 133 375
rect 167 348 179 382
rect 19 249 89 325
rect 19 215 33 249
rect 67 215 89 249
rect 19 195 89 215
rect 133 264 179 348
rect 133 230 145 264
rect 133 161 179 230
rect 35 127 179 161
rect 223 375 224 409
rect 258 375 269 409
rect 223 178 269 375
rect 223 144 231 178
rect 265 144 269 178
rect 35 119 69 127
rect 223 119 269 144
rect 35 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 257 85 269 119
rect 223 69 269 85
rect 307 452 362 489
rect 307 418 328 452
rect 396 483 472 527
rect 822 483 856 527
rect 396 449 422 483
rect 456 449 472 483
rect 579 449 620 483
rect 654 449 778 483
rect 307 415 362 418
rect 307 372 708 415
rect 307 89 341 372
rect 376 321 443 337
rect 376 287 388 321
rect 422 287 443 321
rect 376 157 443 287
rect 477 225 511 372
rect 549 321 630 337
rect 549 287 565 321
rect 599 287 630 321
rect 549 271 630 287
rect 666 321 708 372
rect 744 399 778 449
rect 822 433 856 449
rect 913 472 960 488
rect 1280 485 1314 527
rect 913 438 926 472
rect 1009 438 1035 472
rect 1069 438 1246 472
rect 913 413 960 438
rect 913 399 947 413
rect 744 365 947 399
rect 1077 382 1175 402
rect 666 287 674 321
rect 666 271 708 287
rect 745 288 819 331
rect 745 254 777 288
rect 811 254 819 288
rect 477 191 493 225
rect 527 191 543 225
rect 667 207 701 223
rect 745 207 819 254
rect 913 173 947 365
rect 667 157 701 173
rect 376 123 701 157
rect 745 139 947 173
rect 981 365 1039 381
rect 1015 331 1039 365
rect 1077 365 1133 382
rect 1077 331 1093 365
rect 1127 348 1133 365
rect 1167 348 1175 382
rect 1127 331 1175 348
rect 981 207 1039 331
rect 1209 315 1246 438
rect 1280 417 1314 451
rect 1280 367 1314 383
rect 1371 477 1412 493
rect 1371 443 1378 477
rect 1693 477 1754 527
rect 1209 299 1337 315
rect 1209 297 1287 299
rect 1141 265 1287 297
rect 1321 265 1337 299
rect 1141 263 1337 265
rect 981 191 1107 207
rect 981 178 1073 191
rect 981 144 1031 178
rect 1065 157 1073 178
rect 1065 144 1107 157
rect 981 141 1107 144
rect 745 89 779 139
rect 913 107 947 139
rect 1141 107 1175 263
rect 1371 219 1412 443
rect 1450 433 1486 467
rect 1520 433 1657 467
rect 1446 382 1494 393
rect 1446 348 1448 382
rect 1482 348 1494 382
rect 1446 299 1494 348
rect 1480 265 1494 299
rect 1446 249 1494 265
rect 1547 365 1589 381
rect 1547 331 1548 365
rect 1582 331 1589 365
rect 1209 203 1412 219
rect 1547 207 1589 331
rect 1243 169 1412 203
rect 1209 153 1412 169
rect 103 17 179 59
rect 307 55 331 89
rect 365 55 381 89
rect 415 55 431 89
rect 465 55 481 89
rect 614 55 636 89
rect 670 55 779 89
rect 823 89 863 105
rect 857 55 863 89
rect 913 73 933 107
rect 967 73 983 107
rect 1027 73 1043 107
rect 1077 73 1175 107
rect 1245 101 1319 117
rect 415 17 481 55
rect 823 17 863 55
rect 1245 67 1279 101
rect 1313 67 1319 101
rect 1355 107 1412 153
rect 1450 191 1589 207
rect 1450 157 1456 191
rect 1490 178 1589 191
rect 1450 144 1462 157
rect 1496 144 1589 178
rect 1450 141 1589 144
rect 1623 265 1657 433
rect 1693 443 1719 477
rect 1753 443 1754 477
rect 1693 427 1754 443
rect 1824 475 1881 491
rect 1858 441 1881 475
rect 1824 407 1881 441
rect 1691 373 1824 381
rect 1858 373 1881 407
rect 1691 365 1881 373
rect 1725 331 1881 365
rect 1691 315 1881 331
rect 1918 455 1952 527
rect 1918 375 1952 421
rect 1918 325 1952 341
rect 1986 445 2012 479
rect 2046 445 2094 479
rect 1986 411 2094 445
rect 1986 377 2012 411
rect 2046 377 2094 411
rect 1986 343 2094 377
rect 1844 265 1881 315
rect 1986 309 2012 343
rect 1623 249 1810 265
rect 1623 215 1776 249
rect 1623 199 1810 215
rect 1844 249 2006 265
rect 1844 215 1972 249
rect 1844 199 2006 215
rect 1623 107 1657 199
rect 1844 165 1880 199
rect 1808 162 1880 165
rect 1808 128 1824 162
rect 1858 128 1880 162
rect 1355 73 1402 107
rect 1436 73 1452 107
rect 1491 73 1507 107
rect 1541 73 1657 107
rect 1691 107 1754 123
rect 1691 73 1720 107
rect 1245 17 1319 67
rect 1691 17 1754 73
rect 1808 94 1880 128
rect 1808 60 1824 94
rect 1858 60 1880 94
rect 1918 123 1952 139
rect 1918 17 1952 89
rect 1986 130 2012 164
rect 2046 130 2094 343
rect 1986 96 2094 130
rect 1986 62 2012 96
rect 2046 62 2094 96
rect 1986 61 2094 62
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 133 348 167 382
rect 231 144 265 178
rect 1133 348 1167 382
rect 1031 144 1065 178
rect 1448 348 1482 382
rect 1462 157 1490 178
rect 1490 157 1496 178
rect 1462 144 1496 157
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 121 382 1494 388
rect 121 348 133 382
rect 167 360 1133 382
rect 167 348 179 360
rect 121 342 179 348
rect 1111 348 1133 360
rect 1167 360 1448 382
rect 1167 348 1179 360
rect 1111 342 1179 348
rect 1426 348 1448 360
rect 1482 348 1494 382
rect 1426 342 1494 348
rect 219 178 1508 184
rect 219 144 231 178
rect 265 156 1031 178
rect 265 144 277 156
rect 219 138 277 144
rect 1009 144 1031 156
rect 1065 156 1462 178
rect 1065 144 1077 156
rect 1009 138 1077 144
rect 1446 144 1462 156
rect 1496 144 1508 178
rect 1446 138 1508 144
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfxtp_1
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew signal input
flabel locali s 2046 353 2080 387 0 FreeSans 300 0 0 0 Q
port 9 nsew signal output
flabel locali s 764 221 798 255 0 FreeSans 300 0 0 0 SCD
port 3 nsew signal input
flabel locali s 581 289 615 323 0 FreeSans 300 0 0 0 D
port 2 nsew signal input
flabel locali s 397 152 431 186 0 FreeSans 300 0 0 0 SCE
port 4 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
<< properties >>
string FIXED_BBOX 0 0 2116 544
string GDS_END 2643124
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 2627994
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
