magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 609 157 907 203
rect 1 21 907 157
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 131
rect 287 47 317 131
rect 369 47 399 131
rect 489 47 519 131
rect 588 47 618 131
rect 698 47 728 177
rect 799 47 829 177
<< scpmoshvt >>
rect 81 413 117 497
rect 175 413 211 497
rect 371 413 407 497
rect 481 413 517 497
rect 580 413 616 497
rect 690 297 726 497
rect 791 297 827 497
<< ndiff >>
rect 635 131 698 177
rect 27 93 89 131
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 101 171 131
rect 119 67 129 101
rect 163 67 171 101
rect 119 47 171 67
rect 235 101 287 131
rect 235 67 243 101
rect 277 67 287 101
rect 235 47 287 67
rect 317 47 369 131
rect 399 47 489 131
rect 519 47 588 131
rect 618 93 698 131
rect 618 59 628 93
rect 662 59 698 93
rect 618 47 698 59
rect 728 101 799 177
rect 728 67 745 101
rect 779 67 799 101
rect 728 47 799 67
rect 829 93 881 177
rect 829 59 839 93
rect 873 59 881 93
rect 829 47 881 59
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 413 81 443
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 413 175 451
rect 211 477 371 497
rect 211 443 223 477
rect 257 443 371 477
rect 211 413 371 443
rect 407 485 481 497
rect 407 451 435 485
rect 469 451 481 485
rect 407 413 481 451
rect 517 477 580 497
rect 517 443 534 477
rect 568 443 580 477
rect 517 413 580 443
rect 616 485 690 497
rect 616 451 644 485
rect 678 451 690 485
rect 616 413 690 451
rect 637 297 690 413
rect 726 477 791 497
rect 726 443 745 477
rect 779 443 791 477
rect 726 409 791 443
rect 726 375 745 409
rect 779 375 791 409
rect 726 297 791 375
rect 827 485 881 497
rect 827 451 839 485
rect 873 451 881 485
rect 827 417 881 451
rect 827 383 839 417
rect 873 383 881 417
rect 827 297 881 383
<< ndiffc >>
rect 35 59 69 93
rect 129 67 163 101
rect 243 67 277 101
rect 628 59 662 93
rect 745 67 779 101
rect 839 59 873 93
<< pdiffc >>
rect 35 443 69 477
rect 129 451 163 485
rect 223 443 257 477
rect 435 451 469 485
rect 534 443 568 477
rect 644 451 678 485
rect 745 443 779 477
rect 745 375 779 409
rect 839 451 873 485
rect 839 383 873 417
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 371 497 407 523
rect 481 497 517 523
rect 580 497 616 523
rect 690 497 726 523
rect 791 497 827 523
rect 81 398 117 413
rect 175 398 211 413
rect 371 398 407 413
rect 481 398 517 413
rect 580 398 616 413
rect 79 265 119 398
rect 173 265 213 398
rect 369 349 409 398
rect 369 333 423 349
rect 369 299 379 333
rect 413 299 423 333
rect 369 265 423 299
rect 479 265 519 398
rect 578 265 618 398
rect 690 282 726 297
rect 791 282 827 297
rect 688 265 728 282
rect 789 265 829 282
rect 22 249 119 265
rect 22 215 32 249
rect 66 215 119 249
rect 22 199 119 215
rect 161 249 225 265
rect 161 215 171 249
rect 205 215 225 249
rect 161 199 225 215
rect 89 131 119 199
rect 185 176 225 199
rect 369 231 379 265
rect 413 231 423 265
rect 369 215 423 231
rect 465 249 519 265
rect 465 215 475 249
rect 509 215 519 249
rect 185 146 317 176
rect 287 131 317 146
rect 369 131 399 215
rect 465 199 519 215
rect 564 249 618 265
rect 564 215 574 249
rect 608 215 618 249
rect 564 199 618 215
rect 667 249 829 265
rect 667 215 677 249
rect 711 215 829 249
rect 667 199 829 215
rect 489 131 519 199
rect 588 131 618 199
rect 698 177 728 199
rect 799 177 829 199
rect 89 21 119 47
rect 287 21 317 47
rect 369 21 399 47
rect 489 21 519 47
rect 588 21 618 47
rect 698 21 728 47
rect 799 21 829 47
<< polycont >>
rect 379 299 413 333
rect 32 215 66 249
rect 171 215 205 249
rect 379 231 413 265
rect 475 215 509 249
rect 574 215 608 249
rect 677 215 711 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 35 477 69 493
rect 35 400 69 443
rect 103 485 179 527
rect 103 451 129 485
rect 163 451 179 485
rect 103 439 179 451
rect 223 477 257 493
rect 341 485 485 527
rect 341 451 435 485
rect 469 451 485 485
rect 534 477 572 493
rect 223 417 257 443
rect 568 443 572 477
rect 534 417 572 443
rect 628 485 694 527
rect 628 451 644 485
rect 678 451 694 485
rect 628 439 694 451
rect 738 477 799 493
rect 738 443 745 477
rect 779 443 799 477
rect 35 366 171 400
rect 27 249 67 326
rect 27 215 32 249
rect 66 215 67 249
rect 27 148 67 215
rect 137 265 171 366
rect 223 393 572 417
rect 738 409 799 443
rect 223 383 693 393
rect 223 332 283 383
rect 538 359 693 383
rect 137 249 215 265
rect 137 215 171 249
rect 205 215 215 249
rect 137 199 215 215
rect 137 117 171 199
rect 249 117 283 332
rect 129 101 171 117
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 163 67 171 101
rect 129 51 171 67
rect 239 101 283 117
rect 239 67 243 101
rect 277 67 283 101
rect 379 333 431 349
rect 413 299 431 333
rect 379 265 431 299
rect 413 231 431 265
rect 379 84 431 231
rect 475 249 523 323
rect 509 215 523 249
rect 475 84 523 215
rect 557 249 623 323
rect 557 215 574 249
rect 608 215 623 249
rect 557 129 623 215
rect 659 265 693 359
rect 738 375 745 409
rect 779 375 799 409
rect 738 333 799 375
rect 839 485 890 527
rect 873 451 890 485
rect 839 417 890 451
rect 873 383 890 417
rect 839 367 890 383
rect 738 307 891 333
rect 659 249 711 265
rect 659 215 677 249
rect 659 199 711 215
rect 755 165 891 307
rect 712 128 891 165
rect 712 101 779 128
rect 239 51 283 67
rect 602 59 628 93
rect 662 59 678 93
rect 602 17 678 59
rect 712 67 745 101
rect 712 51 779 67
rect 813 59 839 93
rect 873 59 890 93
rect 813 17 890 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 781 170 781 170 0 FreeSans 200 0 0 0 X
flabel locali s 781 238 781 238 0 FreeSans 200 0 0 0 X
flabel locali s 781 306 781 306 0 FreeSans 200 0 0 0 X
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 742 85 776 119 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 742 357 776 391 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 742 425 776 459 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 558 289 592 323 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 475 84 523 323 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 483 170 483 170 0 FreeSans 200 0 0 0 C
flabel locali s 388 85 422 119 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 388 153 422 187 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 388 221 422 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 388 289 422 323 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 30 153 64 187 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4b_2
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 866268
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 857784
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
