magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 3258 582
<< pwell >>
rect 1 21 3217 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 173 47 203 177
rect 277 47 307 177
rect 361 47 391 177
rect 465 47 495 177
rect 549 47 579 177
rect 653 47 683 177
rect 737 47 767 177
rect 841 47 871 177
rect 925 47 955 177
rect 1029 47 1059 177
rect 1113 47 1143 177
rect 1217 47 1247 177
rect 1301 47 1331 177
rect 1405 47 1435 177
rect 1489 47 1519 177
rect 1697 47 1727 177
rect 1781 47 1811 177
rect 1885 47 1915 177
rect 1969 47 1999 177
rect 2073 47 2103 177
rect 2157 47 2187 177
rect 2261 47 2291 177
rect 2345 47 2375 177
rect 2449 47 2479 177
rect 2533 47 2563 177
rect 2637 47 2667 177
rect 2721 47 2751 177
rect 2825 47 2855 177
rect 2909 47 2939 177
rect 3013 47 3043 177
rect 3097 47 3127 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
rect 1209 297 1245 497
rect 1303 297 1339 497
rect 1397 297 1433 497
rect 1491 297 1527 497
rect 1689 297 1725 497
rect 1783 297 1819 497
rect 1877 297 1913 497
rect 1971 297 2007 497
rect 2065 297 2101 497
rect 2159 297 2195 497
rect 2253 297 2289 497
rect 2347 297 2383 497
rect 2441 297 2477 497
rect 2535 297 2571 497
rect 2629 297 2665 497
rect 2723 297 2759 497
rect 2817 297 2853 497
rect 2911 297 2947 497
rect 3005 297 3041 497
rect 3099 297 3135 497
<< ndiff >>
rect 27 163 89 177
rect 27 129 35 163
rect 69 129 89 163
rect 27 95 89 129
rect 27 61 35 95
rect 69 61 89 95
rect 27 47 89 61
rect 119 163 173 177
rect 119 129 129 163
rect 163 129 173 163
rect 119 95 173 129
rect 119 61 129 95
rect 163 61 173 95
rect 119 47 173 61
rect 203 95 277 177
rect 203 61 223 95
rect 257 61 277 95
rect 203 47 277 61
rect 307 163 361 177
rect 307 129 317 163
rect 351 129 361 163
rect 307 95 361 129
rect 307 61 317 95
rect 351 61 361 95
rect 307 47 361 61
rect 391 95 465 177
rect 391 61 411 95
rect 445 61 465 95
rect 391 47 465 61
rect 495 163 549 177
rect 495 129 505 163
rect 539 129 549 163
rect 495 95 549 129
rect 495 61 505 95
rect 539 61 549 95
rect 495 47 549 61
rect 579 95 653 177
rect 579 61 599 95
rect 633 61 653 95
rect 579 47 653 61
rect 683 163 737 177
rect 683 129 693 163
rect 727 129 737 163
rect 683 95 737 129
rect 683 61 693 95
rect 727 61 737 95
rect 683 47 737 61
rect 767 95 841 177
rect 767 61 787 95
rect 821 61 841 95
rect 767 47 841 61
rect 871 163 925 177
rect 871 129 881 163
rect 915 129 925 163
rect 871 95 925 129
rect 871 61 881 95
rect 915 61 925 95
rect 871 47 925 61
rect 955 95 1029 177
rect 955 61 975 95
rect 1009 61 1029 95
rect 955 47 1029 61
rect 1059 163 1113 177
rect 1059 129 1069 163
rect 1103 129 1113 163
rect 1059 95 1113 129
rect 1059 61 1069 95
rect 1103 61 1113 95
rect 1059 47 1113 61
rect 1143 95 1217 177
rect 1143 61 1163 95
rect 1197 61 1217 95
rect 1143 47 1217 61
rect 1247 163 1301 177
rect 1247 129 1257 163
rect 1291 129 1301 163
rect 1247 95 1301 129
rect 1247 61 1257 95
rect 1291 61 1301 95
rect 1247 47 1301 61
rect 1331 95 1405 177
rect 1331 61 1351 95
rect 1385 61 1405 95
rect 1331 47 1405 61
rect 1435 163 1489 177
rect 1435 129 1445 163
rect 1479 129 1489 163
rect 1435 95 1489 129
rect 1435 61 1445 95
rect 1479 61 1489 95
rect 1435 47 1489 61
rect 1519 95 1697 177
rect 1519 61 1539 95
rect 1573 61 1643 95
rect 1677 61 1697 95
rect 1519 47 1697 61
rect 1727 163 1781 177
rect 1727 129 1737 163
rect 1771 129 1781 163
rect 1727 95 1781 129
rect 1727 61 1737 95
rect 1771 61 1781 95
rect 1727 47 1781 61
rect 1811 95 1885 177
rect 1811 61 1831 95
rect 1865 61 1885 95
rect 1811 47 1885 61
rect 1915 163 1969 177
rect 1915 129 1925 163
rect 1959 129 1969 163
rect 1915 95 1969 129
rect 1915 61 1925 95
rect 1959 61 1969 95
rect 1915 47 1969 61
rect 1999 95 2073 177
rect 1999 61 2019 95
rect 2053 61 2073 95
rect 1999 47 2073 61
rect 2103 163 2157 177
rect 2103 129 2113 163
rect 2147 129 2157 163
rect 2103 95 2157 129
rect 2103 61 2113 95
rect 2147 61 2157 95
rect 2103 47 2157 61
rect 2187 95 2261 177
rect 2187 61 2207 95
rect 2241 61 2261 95
rect 2187 47 2261 61
rect 2291 163 2345 177
rect 2291 129 2301 163
rect 2335 129 2345 163
rect 2291 95 2345 129
rect 2291 61 2301 95
rect 2335 61 2345 95
rect 2291 47 2345 61
rect 2375 95 2449 177
rect 2375 61 2395 95
rect 2429 61 2449 95
rect 2375 47 2449 61
rect 2479 163 2533 177
rect 2479 129 2489 163
rect 2523 129 2533 163
rect 2479 95 2533 129
rect 2479 61 2489 95
rect 2523 61 2533 95
rect 2479 47 2533 61
rect 2563 95 2637 177
rect 2563 61 2583 95
rect 2617 61 2637 95
rect 2563 47 2637 61
rect 2667 163 2721 177
rect 2667 129 2677 163
rect 2711 129 2721 163
rect 2667 95 2721 129
rect 2667 61 2677 95
rect 2711 61 2721 95
rect 2667 47 2721 61
rect 2751 95 2825 177
rect 2751 61 2771 95
rect 2805 61 2825 95
rect 2751 47 2825 61
rect 2855 163 2909 177
rect 2855 129 2865 163
rect 2899 129 2909 163
rect 2855 95 2909 129
rect 2855 61 2865 95
rect 2899 61 2909 95
rect 2855 47 2909 61
rect 2939 95 3013 177
rect 2939 61 2961 95
rect 2995 61 3013 95
rect 2939 47 3013 61
rect 3043 163 3097 177
rect 3043 129 3053 163
rect 3087 129 3097 163
rect 3043 95 3097 129
rect 3043 61 3053 95
rect 3087 61 3097 95
rect 3043 47 3097 61
rect 3127 163 3191 177
rect 3127 129 3149 163
rect 3183 129 3191 163
rect 3127 95 3191 129
rect 3127 61 3149 95
rect 3183 61 3191 95
rect 3127 47 3191 61
<< pdiff >>
rect 27 479 81 497
rect 27 445 35 479
rect 69 445 81 479
rect 27 411 81 445
rect 27 377 35 411
rect 69 377 81 411
rect 27 343 81 377
rect 27 309 35 343
rect 69 309 81 343
rect 27 297 81 309
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 297 175 375
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 409 269 443
rect 211 375 223 409
rect 257 375 269 409
rect 211 341 269 375
rect 211 307 223 341
rect 257 307 269 341
rect 211 297 269 307
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 409 363 443
rect 305 375 317 409
rect 351 375 363 409
rect 305 297 363 375
rect 399 477 457 497
rect 399 443 411 477
rect 445 443 457 477
rect 399 409 457 443
rect 399 375 411 409
rect 445 375 457 409
rect 399 341 457 375
rect 399 307 411 341
rect 445 307 457 341
rect 399 297 457 307
rect 493 477 551 497
rect 493 443 505 477
rect 539 443 551 477
rect 493 409 551 443
rect 493 375 505 409
rect 539 375 551 409
rect 493 297 551 375
rect 587 477 645 497
rect 587 443 599 477
rect 633 443 645 477
rect 587 409 645 443
rect 587 375 599 409
rect 633 375 645 409
rect 587 341 645 375
rect 587 307 599 341
rect 633 307 645 341
rect 587 297 645 307
rect 681 477 739 497
rect 681 443 693 477
rect 727 443 739 477
rect 681 409 739 443
rect 681 375 693 409
rect 727 375 739 409
rect 681 297 739 375
rect 775 477 833 497
rect 775 443 787 477
rect 821 443 833 477
rect 775 409 833 443
rect 775 375 787 409
rect 821 375 833 409
rect 775 341 833 375
rect 775 307 787 341
rect 821 307 833 341
rect 775 297 833 307
rect 869 409 927 497
rect 869 375 881 409
rect 915 375 927 409
rect 869 341 927 375
rect 869 307 881 341
rect 915 307 927 341
rect 869 297 927 307
rect 963 477 1021 497
rect 963 443 975 477
rect 1009 443 1021 477
rect 963 409 1021 443
rect 963 375 975 409
rect 1009 375 1021 409
rect 963 297 1021 375
rect 1057 409 1115 497
rect 1057 375 1069 409
rect 1103 375 1115 409
rect 1057 341 1115 375
rect 1057 307 1069 341
rect 1103 307 1115 341
rect 1057 297 1115 307
rect 1151 477 1209 497
rect 1151 443 1163 477
rect 1197 443 1209 477
rect 1151 409 1209 443
rect 1151 375 1163 409
rect 1197 375 1209 409
rect 1151 297 1209 375
rect 1245 409 1303 497
rect 1245 375 1257 409
rect 1291 375 1303 409
rect 1245 341 1303 375
rect 1245 307 1257 341
rect 1291 307 1303 341
rect 1245 297 1303 307
rect 1339 477 1397 497
rect 1339 443 1351 477
rect 1385 443 1397 477
rect 1339 409 1397 443
rect 1339 375 1351 409
rect 1385 375 1397 409
rect 1339 297 1397 375
rect 1433 409 1491 497
rect 1433 375 1445 409
rect 1479 375 1491 409
rect 1433 341 1491 375
rect 1433 307 1445 341
rect 1479 307 1491 341
rect 1433 297 1491 307
rect 1527 477 1581 497
rect 1527 443 1539 477
rect 1573 443 1581 477
rect 1527 409 1581 443
rect 1527 375 1539 409
rect 1573 375 1581 409
rect 1527 297 1581 375
rect 1635 477 1689 497
rect 1635 443 1643 477
rect 1677 443 1689 477
rect 1635 409 1689 443
rect 1635 375 1643 409
rect 1677 375 1689 409
rect 1635 297 1689 375
rect 1725 409 1783 497
rect 1725 375 1737 409
rect 1771 375 1783 409
rect 1725 341 1783 375
rect 1725 307 1737 341
rect 1771 307 1783 341
rect 1725 297 1783 307
rect 1819 477 1877 497
rect 1819 443 1831 477
rect 1865 443 1877 477
rect 1819 409 1877 443
rect 1819 375 1831 409
rect 1865 375 1877 409
rect 1819 297 1877 375
rect 1913 409 1971 497
rect 1913 375 1925 409
rect 1959 375 1971 409
rect 1913 341 1971 375
rect 1913 307 1925 341
rect 1959 307 1971 341
rect 1913 297 1971 307
rect 2007 477 2065 497
rect 2007 443 2019 477
rect 2053 443 2065 477
rect 2007 409 2065 443
rect 2007 375 2019 409
rect 2053 375 2065 409
rect 2007 297 2065 375
rect 2101 409 2159 497
rect 2101 375 2113 409
rect 2147 375 2159 409
rect 2101 341 2159 375
rect 2101 307 2113 341
rect 2147 307 2159 341
rect 2101 297 2159 307
rect 2195 477 2253 497
rect 2195 443 2207 477
rect 2241 443 2253 477
rect 2195 409 2253 443
rect 2195 375 2207 409
rect 2241 375 2253 409
rect 2195 297 2253 375
rect 2289 409 2347 497
rect 2289 375 2301 409
rect 2335 375 2347 409
rect 2289 341 2347 375
rect 2289 307 2301 341
rect 2335 307 2347 341
rect 2289 297 2347 307
rect 2383 477 2441 497
rect 2383 443 2395 477
rect 2429 443 2441 477
rect 2383 409 2441 443
rect 2383 375 2395 409
rect 2429 375 2441 409
rect 2383 341 2441 375
rect 2383 307 2395 341
rect 2429 307 2441 341
rect 2383 297 2441 307
rect 2477 409 2535 497
rect 2477 375 2489 409
rect 2523 375 2535 409
rect 2477 341 2535 375
rect 2477 307 2489 341
rect 2523 307 2535 341
rect 2477 297 2535 307
rect 2571 477 2629 497
rect 2571 443 2583 477
rect 2617 443 2629 477
rect 2571 409 2629 443
rect 2571 375 2583 409
rect 2617 375 2629 409
rect 2571 297 2629 375
rect 2665 409 2723 497
rect 2665 375 2677 409
rect 2711 375 2723 409
rect 2665 341 2723 375
rect 2665 307 2677 341
rect 2711 307 2723 341
rect 2665 297 2723 307
rect 2759 477 2817 497
rect 2759 443 2771 477
rect 2805 443 2817 477
rect 2759 409 2817 443
rect 2759 375 2771 409
rect 2805 375 2817 409
rect 2759 297 2817 375
rect 2853 409 2911 497
rect 2853 375 2865 409
rect 2899 375 2911 409
rect 2853 341 2911 375
rect 2853 307 2865 341
rect 2899 307 2911 341
rect 2853 297 2911 307
rect 2947 477 3005 497
rect 2947 443 2961 477
rect 2995 443 3005 477
rect 2947 409 3005 443
rect 2947 375 2961 409
rect 2995 375 3005 409
rect 2947 297 3005 375
rect 3041 409 3099 497
rect 3041 375 3053 409
rect 3087 375 3099 409
rect 3041 341 3099 375
rect 3041 307 3053 341
rect 3087 307 3099 341
rect 3041 297 3099 307
rect 3135 479 3191 497
rect 3135 445 3149 479
rect 3183 445 3191 479
rect 3135 411 3191 445
rect 3135 377 3149 411
rect 3183 377 3191 411
rect 3135 343 3191 377
rect 3135 309 3149 343
rect 3183 309 3191 343
rect 3135 297 3191 309
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 129 129 163 163
rect 129 61 163 95
rect 223 61 257 95
rect 317 129 351 163
rect 317 61 351 95
rect 411 61 445 95
rect 505 129 539 163
rect 505 61 539 95
rect 599 61 633 95
rect 693 129 727 163
rect 693 61 727 95
rect 787 61 821 95
rect 881 129 915 163
rect 881 61 915 95
rect 975 61 1009 95
rect 1069 129 1103 163
rect 1069 61 1103 95
rect 1163 61 1197 95
rect 1257 129 1291 163
rect 1257 61 1291 95
rect 1351 61 1385 95
rect 1445 129 1479 163
rect 1445 61 1479 95
rect 1539 61 1573 95
rect 1643 61 1677 95
rect 1737 129 1771 163
rect 1737 61 1771 95
rect 1831 61 1865 95
rect 1925 129 1959 163
rect 1925 61 1959 95
rect 2019 61 2053 95
rect 2113 129 2147 163
rect 2113 61 2147 95
rect 2207 61 2241 95
rect 2301 129 2335 163
rect 2301 61 2335 95
rect 2395 61 2429 95
rect 2489 129 2523 163
rect 2489 61 2523 95
rect 2583 61 2617 95
rect 2677 129 2711 163
rect 2677 61 2711 95
rect 2771 61 2805 95
rect 2865 129 2899 163
rect 2865 61 2899 95
rect 2961 61 2995 95
rect 3053 129 3087 163
rect 3053 61 3087 95
rect 3149 129 3183 163
rect 3149 61 3183 95
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 129 443 163 477
rect 129 375 163 409
rect 223 443 257 477
rect 223 375 257 409
rect 223 307 257 341
rect 317 443 351 477
rect 317 375 351 409
rect 411 443 445 477
rect 411 375 445 409
rect 411 307 445 341
rect 505 443 539 477
rect 505 375 539 409
rect 599 443 633 477
rect 599 375 633 409
rect 599 307 633 341
rect 693 443 727 477
rect 693 375 727 409
rect 787 443 821 477
rect 787 375 821 409
rect 787 307 821 341
rect 881 375 915 409
rect 881 307 915 341
rect 975 443 1009 477
rect 975 375 1009 409
rect 1069 375 1103 409
rect 1069 307 1103 341
rect 1163 443 1197 477
rect 1163 375 1197 409
rect 1257 375 1291 409
rect 1257 307 1291 341
rect 1351 443 1385 477
rect 1351 375 1385 409
rect 1445 375 1479 409
rect 1445 307 1479 341
rect 1539 443 1573 477
rect 1539 375 1573 409
rect 1643 443 1677 477
rect 1643 375 1677 409
rect 1737 375 1771 409
rect 1737 307 1771 341
rect 1831 443 1865 477
rect 1831 375 1865 409
rect 1925 375 1959 409
rect 1925 307 1959 341
rect 2019 443 2053 477
rect 2019 375 2053 409
rect 2113 375 2147 409
rect 2113 307 2147 341
rect 2207 443 2241 477
rect 2207 375 2241 409
rect 2301 375 2335 409
rect 2301 307 2335 341
rect 2395 443 2429 477
rect 2395 375 2429 409
rect 2395 307 2429 341
rect 2489 375 2523 409
rect 2489 307 2523 341
rect 2583 443 2617 477
rect 2583 375 2617 409
rect 2677 375 2711 409
rect 2677 307 2711 341
rect 2771 443 2805 477
rect 2771 375 2805 409
rect 2865 375 2899 409
rect 2865 307 2899 341
rect 2961 443 2995 477
rect 2961 375 2995 409
rect 3053 375 3087 409
rect 3053 307 3087 341
rect 3149 445 3183 479
rect 3149 377 3183 411
rect 3149 309 3183 343
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 1209 497 1245 523
rect 1303 497 1339 523
rect 1397 497 1433 523
rect 1491 497 1527 523
rect 1689 497 1725 523
rect 1783 497 1819 523
rect 1877 497 1913 523
rect 1971 497 2007 523
rect 2065 497 2101 523
rect 2159 497 2195 523
rect 2253 497 2289 523
rect 2347 497 2383 523
rect 2441 497 2477 523
rect 2535 497 2571 523
rect 2629 497 2665 523
rect 2723 497 2759 523
rect 2817 497 2853 523
rect 2911 497 2947 523
rect 3005 497 3041 523
rect 3099 497 3135 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 1209 282 1245 297
rect 1303 282 1339 297
rect 1397 282 1433 297
rect 1491 282 1527 297
rect 1689 282 1725 297
rect 1783 282 1819 297
rect 1877 282 1913 297
rect 1971 282 2007 297
rect 2065 282 2101 297
rect 2159 282 2195 297
rect 2253 282 2289 297
rect 2347 282 2383 297
rect 2441 282 2477 297
rect 2535 282 2571 297
rect 2629 282 2665 297
rect 2723 282 2759 297
rect 2817 282 2853 297
rect 2911 282 2947 297
rect 3005 282 3041 297
rect 3099 282 3135 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 79 249 777 265
rect 79 215 97 249
rect 131 215 165 249
rect 199 215 233 249
rect 267 215 301 249
rect 335 215 369 249
rect 403 215 437 249
rect 471 215 505 249
rect 539 215 573 249
rect 607 215 641 249
rect 675 215 709 249
rect 743 215 777 249
rect 79 199 777 215
rect 831 265 871 282
rect 925 265 965 282
rect 1019 265 1059 282
rect 1113 265 1153 282
rect 1207 265 1247 282
rect 1301 265 1341 282
rect 1395 265 1435 282
rect 1489 265 1529 282
rect 831 249 1529 265
rect 831 215 865 249
rect 899 215 933 249
rect 967 215 1001 249
rect 1035 215 1069 249
rect 1103 215 1137 249
rect 1171 215 1205 249
rect 1239 215 1273 249
rect 1307 215 1341 249
rect 1375 215 1409 249
rect 1443 215 1477 249
rect 1511 215 1529 249
rect 831 199 1529 215
rect 1687 265 1727 282
rect 1781 265 1821 282
rect 1875 265 1915 282
rect 1969 265 2009 282
rect 2063 265 2103 282
rect 2157 265 2197 282
rect 2251 265 2291 282
rect 2345 265 2385 282
rect 1687 249 2385 265
rect 1687 215 1705 249
rect 1739 215 1773 249
rect 1807 215 1841 249
rect 1875 215 1909 249
rect 1943 215 1977 249
rect 2011 215 2045 249
rect 2079 215 2113 249
rect 2147 215 2181 249
rect 2215 215 2249 249
rect 2283 215 2317 249
rect 2351 215 2385 249
rect 1687 199 2385 215
rect 2439 265 2479 282
rect 2533 265 2573 282
rect 2627 265 2667 282
rect 2721 265 2761 282
rect 2815 265 2855 282
rect 2909 265 2949 282
rect 3003 265 3043 282
rect 3097 265 3137 282
rect 2439 249 3137 265
rect 2439 215 2613 249
rect 2647 215 2681 249
rect 2715 215 2749 249
rect 2783 215 2817 249
rect 2851 215 2885 249
rect 2919 215 2953 249
rect 2987 215 3021 249
rect 3055 215 3137 249
rect 2439 199 3137 215
rect 89 177 119 199
rect 173 177 203 199
rect 277 177 307 199
rect 361 177 391 199
rect 465 177 495 199
rect 549 177 579 199
rect 653 177 683 199
rect 737 177 767 199
rect 841 177 871 199
rect 925 177 955 199
rect 1029 177 1059 199
rect 1113 177 1143 199
rect 1217 177 1247 199
rect 1301 177 1331 199
rect 1405 177 1435 199
rect 1489 177 1519 199
rect 1697 177 1727 199
rect 1781 177 1811 199
rect 1885 177 1915 199
rect 1969 177 1999 199
rect 2073 177 2103 199
rect 2157 177 2187 199
rect 2261 177 2291 199
rect 2345 177 2375 199
rect 2449 177 2479 199
rect 2533 177 2563 199
rect 2637 177 2667 199
rect 2721 177 2751 199
rect 2825 177 2855 199
rect 2909 177 2939 199
rect 3013 177 3043 199
rect 3097 177 3127 199
rect 89 21 119 47
rect 173 21 203 47
rect 277 21 307 47
rect 361 21 391 47
rect 465 21 495 47
rect 549 21 579 47
rect 653 21 683 47
rect 737 21 767 47
rect 841 21 871 47
rect 925 21 955 47
rect 1029 21 1059 47
rect 1113 21 1143 47
rect 1217 21 1247 47
rect 1301 21 1331 47
rect 1405 21 1435 47
rect 1489 21 1519 47
rect 1697 21 1727 47
rect 1781 21 1811 47
rect 1885 21 1915 47
rect 1969 21 1999 47
rect 2073 21 2103 47
rect 2157 21 2187 47
rect 2261 21 2291 47
rect 2345 21 2375 47
rect 2449 21 2479 47
rect 2533 21 2563 47
rect 2637 21 2667 47
rect 2721 21 2751 47
rect 2825 21 2855 47
rect 2909 21 2939 47
rect 3013 21 3043 47
rect 3097 21 3127 47
<< polycont >>
rect 97 215 131 249
rect 165 215 199 249
rect 233 215 267 249
rect 301 215 335 249
rect 369 215 403 249
rect 437 215 471 249
rect 505 215 539 249
rect 573 215 607 249
rect 641 215 675 249
rect 709 215 743 249
rect 865 215 899 249
rect 933 215 967 249
rect 1001 215 1035 249
rect 1069 215 1103 249
rect 1137 215 1171 249
rect 1205 215 1239 249
rect 1273 215 1307 249
rect 1341 215 1375 249
rect 1409 215 1443 249
rect 1477 215 1511 249
rect 1705 215 1739 249
rect 1773 215 1807 249
rect 1841 215 1875 249
rect 1909 215 1943 249
rect 1977 215 2011 249
rect 2045 215 2079 249
rect 2113 215 2147 249
rect 2181 215 2215 249
rect 2249 215 2283 249
rect 2317 215 2351 249
rect 2613 215 2647 249
rect 2681 215 2715 249
rect 2749 215 2783 249
rect 2817 215 2851 249
rect 2885 215 2919 249
rect 2953 215 2987 249
rect 3021 215 3055 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3220 561
rect 19 479 85 493
rect 19 445 35 479
rect 69 445 85 479
rect 19 411 85 445
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 121 477 171 527
rect 121 443 129 477
rect 163 443 171 477
rect 121 409 171 443
rect 121 375 129 409
rect 163 375 171 409
rect 121 359 171 375
rect 215 477 265 493
rect 215 443 223 477
rect 257 443 265 477
rect 215 409 265 443
rect 215 375 223 409
rect 257 375 265 409
rect 19 309 35 343
rect 69 325 85 343
rect 215 341 265 375
rect 309 477 359 527
rect 309 443 317 477
rect 351 443 359 477
rect 309 409 359 443
rect 309 375 317 409
rect 351 375 359 409
rect 309 359 359 375
rect 403 477 453 493
rect 403 443 411 477
rect 445 443 453 477
rect 403 409 453 443
rect 403 375 411 409
rect 445 375 453 409
rect 215 325 223 341
rect 69 309 223 325
rect 19 307 223 309
rect 257 325 265 341
rect 403 341 453 375
rect 497 477 547 527
rect 497 443 505 477
rect 539 443 547 477
rect 497 409 547 443
rect 497 375 505 409
rect 539 375 547 409
rect 497 359 547 375
rect 591 477 641 493
rect 591 443 599 477
rect 633 443 641 477
rect 591 409 641 443
rect 591 375 599 409
rect 633 375 641 409
rect 403 325 411 341
rect 257 307 411 325
rect 445 325 453 341
rect 591 341 641 375
rect 685 477 735 527
rect 685 443 693 477
rect 727 443 735 477
rect 685 409 735 443
rect 685 375 693 409
rect 727 375 735 409
rect 685 359 735 375
rect 779 477 1589 493
rect 779 443 787 477
rect 821 459 975 477
rect 821 443 829 459
rect 779 409 829 443
rect 967 443 975 459
rect 1009 459 1163 477
rect 1009 443 1017 459
rect 779 375 787 409
rect 821 375 829 409
rect 591 325 599 341
rect 445 307 599 325
rect 633 325 641 341
rect 779 341 829 375
rect 779 325 787 341
rect 633 307 787 325
rect 821 307 829 341
rect 19 291 829 307
rect 873 409 923 425
rect 873 375 881 409
rect 915 375 923 409
rect 873 341 923 375
rect 967 409 1017 443
rect 1155 443 1163 459
rect 1197 459 1351 477
rect 1197 443 1205 459
rect 967 375 975 409
rect 1009 375 1017 409
rect 967 359 1017 375
rect 1061 409 1111 425
rect 1061 375 1069 409
rect 1103 375 1111 409
rect 873 307 881 341
rect 915 325 923 341
rect 1061 341 1111 375
rect 1155 409 1205 443
rect 1343 443 1351 459
rect 1385 459 1539 477
rect 1385 443 1393 459
rect 1155 375 1163 409
rect 1197 375 1205 409
rect 1155 359 1205 375
rect 1249 409 1299 425
rect 1249 375 1257 409
rect 1291 375 1299 409
rect 1061 325 1069 341
rect 915 307 1069 325
rect 1103 325 1111 341
rect 1249 341 1299 375
rect 1343 409 1393 443
rect 1531 443 1539 459
rect 1573 443 1589 477
rect 1343 375 1351 409
rect 1385 375 1393 409
rect 1343 359 1393 375
rect 1437 409 1487 425
rect 1437 375 1445 409
rect 1479 375 1487 409
rect 1249 325 1257 341
rect 1103 307 1257 325
rect 1291 325 1299 341
rect 1437 341 1487 375
rect 1531 409 1589 443
rect 1531 375 1539 409
rect 1573 375 1589 409
rect 1531 359 1589 375
rect 1627 479 3199 493
rect 1627 477 3149 479
rect 1627 443 1643 477
rect 1677 459 1831 477
rect 1677 443 1685 459
rect 1627 409 1685 443
rect 1815 443 1831 459
rect 1865 459 2019 477
rect 1865 443 1873 459
rect 1627 375 1643 409
rect 1677 375 1685 409
rect 1627 359 1685 375
rect 1729 409 1779 425
rect 1729 375 1737 409
rect 1771 375 1779 409
rect 1437 325 1445 341
rect 1291 307 1445 325
rect 1479 325 1487 341
rect 1729 341 1779 375
rect 1815 409 1873 443
rect 2011 443 2019 459
rect 2053 459 2207 477
rect 2053 443 2061 459
rect 1815 375 1831 409
rect 1865 375 1873 409
rect 1815 359 1873 375
rect 1917 409 1967 425
rect 1917 375 1925 409
rect 1959 375 1967 409
rect 1729 325 1737 341
rect 1479 307 1737 325
rect 1771 325 1779 341
rect 1917 341 1967 375
rect 2011 409 2061 443
rect 2199 443 2207 459
rect 2241 459 2395 477
rect 2241 443 2249 459
rect 2011 375 2019 409
rect 2053 375 2061 409
rect 2011 359 2061 375
rect 2105 409 2155 425
rect 2105 375 2113 409
rect 2147 375 2155 409
rect 1917 325 1925 341
rect 1771 307 1925 325
rect 1959 325 1967 341
rect 2105 341 2155 375
rect 2199 409 2249 443
rect 2387 443 2395 459
rect 2429 459 2583 477
rect 2429 443 2437 459
rect 2199 375 2207 409
rect 2241 375 2249 409
rect 2199 359 2249 375
rect 2293 409 2343 425
rect 2293 375 2301 409
rect 2335 375 2343 409
rect 2105 325 2113 341
rect 1959 307 2113 325
rect 2147 325 2155 341
rect 2293 341 2343 375
rect 2293 325 2301 341
rect 2147 307 2301 325
rect 2335 307 2343 341
rect 873 291 2343 307
rect 2387 409 2437 443
rect 2575 443 2583 459
rect 2617 459 2771 477
rect 2617 443 2625 459
rect 2387 375 2395 409
rect 2429 375 2437 409
rect 2387 341 2437 375
rect 2387 307 2395 341
rect 2429 307 2437 341
rect 2387 291 2437 307
rect 2481 409 2531 425
rect 2481 375 2489 409
rect 2523 375 2531 409
rect 2481 341 2531 375
rect 2575 409 2625 443
rect 2763 443 2771 459
rect 2805 459 2961 477
rect 2805 443 2813 459
rect 2575 375 2583 409
rect 2617 375 2625 409
rect 2575 359 2625 375
rect 2669 409 2719 425
rect 2669 375 2677 409
rect 2711 375 2719 409
rect 2481 307 2489 341
rect 2523 325 2531 341
rect 2669 341 2719 375
rect 2763 409 2813 443
rect 2951 443 2961 459
rect 2995 459 3149 477
rect 2995 443 3001 459
rect 2763 375 2771 409
rect 2805 375 2813 409
rect 2763 359 2813 375
rect 2857 409 2907 425
rect 2857 375 2865 409
rect 2899 375 2907 409
rect 2669 325 2677 341
rect 2523 307 2677 325
rect 2711 325 2719 341
rect 2857 341 2907 375
rect 2951 409 3001 443
rect 3139 445 3149 459
rect 3183 445 3199 479
rect 2951 375 2961 409
rect 2995 375 3001 409
rect 2951 359 3001 375
rect 3045 409 3095 425
rect 3045 375 3053 409
rect 3087 375 3095 409
rect 2857 325 2865 341
rect 2711 307 2865 325
rect 2899 325 2907 341
rect 3045 341 3095 375
rect 3045 325 3053 341
rect 2899 307 3053 325
rect 3087 307 3095 341
rect 2481 291 3095 307
rect 3139 411 3199 445
rect 3139 377 3149 411
rect 3183 377 3199 411
rect 3139 343 3199 377
rect 3139 309 3149 343
rect 3183 309 3199 343
rect 3139 293 3199 309
rect 81 249 759 257
rect 81 215 97 249
rect 131 215 165 249
rect 199 215 233 249
rect 267 215 301 249
rect 335 215 369 249
rect 403 215 437 249
rect 471 215 505 249
rect 539 215 573 249
rect 607 215 641 249
rect 675 215 709 249
rect 743 215 759 249
rect 849 249 1527 257
rect 849 215 865 249
rect 899 215 933 249
rect 967 215 1001 249
rect 1035 215 1069 249
rect 1103 215 1137 249
rect 1171 215 1205 249
rect 1239 215 1273 249
rect 1307 215 1341 249
rect 1375 215 1409 249
rect 1443 215 1477 249
rect 1511 215 1527 249
rect 1689 249 2367 257
rect 1689 215 1705 249
rect 1739 215 1773 249
rect 1807 215 1841 249
rect 1875 215 1909 249
rect 1943 215 1977 249
rect 2011 215 2045 249
rect 2079 215 2113 249
rect 2147 215 2181 249
rect 2215 215 2249 249
rect 2283 215 2317 249
rect 2351 215 2367 249
rect 2481 181 2563 291
rect 2597 249 3071 257
rect 2597 215 2613 249
rect 2647 215 2681 249
rect 2715 215 2749 249
rect 2783 215 2817 249
rect 2851 215 2885 249
rect 2919 215 2953 249
rect 2987 215 3021 249
rect 3055 215 3071 249
rect 27 163 79 181
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 17 79 61
rect 113 163 3103 181
rect 113 129 129 163
rect 163 145 317 163
rect 163 129 179 145
rect 113 95 179 129
rect 301 129 317 145
rect 351 145 505 163
rect 351 129 367 145
rect 113 61 129 95
rect 163 61 179 95
rect 113 51 179 61
rect 213 95 267 111
rect 213 61 223 95
rect 257 61 267 95
rect 213 17 267 61
rect 301 95 367 129
rect 489 129 505 145
rect 539 145 693 163
rect 539 129 555 145
rect 301 61 317 95
rect 351 61 367 95
rect 301 51 367 61
rect 401 95 455 111
rect 401 61 411 95
rect 445 61 455 95
rect 401 17 455 61
rect 489 95 555 129
rect 677 129 693 145
rect 727 145 881 163
rect 727 129 743 145
rect 489 61 505 95
rect 539 61 555 95
rect 489 51 555 61
rect 589 95 643 111
rect 589 61 599 95
rect 633 61 643 95
rect 589 17 643 61
rect 677 95 743 129
rect 865 129 881 145
rect 915 145 1069 163
rect 915 129 931 145
rect 677 61 693 95
rect 727 61 743 95
rect 677 51 743 61
rect 777 95 831 111
rect 777 61 787 95
rect 821 61 831 95
rect 777 17 831 61
rect 865 95 931 129
rect 1053 129 1069 145
rect 1103 145 1257 163
rect 1103 129 1119 145
rect 865 61 881 95
rect 915 61 931 95
rect 865 51 931 61
rect 965 95 1019 111
rect 965 61 975 95
rect 1009 61 1019 95
rect 965 17 1019 61
rect 1053 95 1119 129
rect 1241 129 1257 145
rect 1291 145 1445 163
rect 1291 129 1307 145
rect 1053 61 1069 95
rect 1103 61 1119 95
rect 1053 51 1119 61
rect 1153 95 1207 111
rect 1153 61 1163 95
rect 1197 61 1207 95
rect 1153 17 1207 61
rect 1241 95 1307 129
rect 1429 129 1445 145
rect 1479 145 1737 163
rect 1479 129 1495 145
rect 1241 61 1257 95
rect 1291 61 1307 95
rect 1241 51 1307 61
rect 1341 95 1395 111
rect 1341 61 1351 95
rect 1385 61 1395 95
rect 1341 17 1395 61
rect 1429 95 1495 129
rect 1721 129 1737 145
rect 1771 145 1925 163
rect 1771 129 1787 145
rect 1429 61 1445 95
rect 1479 61 1495 95
rect 1429 51 1495 61
rect 1529 95 1687 111
rect 1529 61 1539 95
rect 1573 61 1643 95
rect 1677 61 1687 95
rect 1529 17 1687 61
rect 1721 95 1787 129
rect 1909 129 1925 145
rect 1959 145 2113 163
rect 1959 129 1975 145
rect 1721 61 1737 95
rect 1771 61 1787 95
rect 1721 51 1787 61
rect 1821 95 1875 111
rect 1821 61 1831 95
rect 1865 61 1875 95
rect 1821 17 1875 61
rect 1909 95 1975 129
rect 2097 129 2113 145
rect 2147 145 2301 163
rect 2147 129 2163 145
rect 1909 61 1925 95
rect 1959 61 1975 95
rect 1909 51 1975 61
rect 2009 95 2063 111
rect 2009 61 2019 95
rect 2053 61 2063 95
rect 2009 17 2063 61
rect 2097 95 2163 129
rect 2285 129 2301 145
rect 2335 145 2489 163
rect 2335 129 2351 145
rect 2097 61 2113 95
rect 2147 61 2163 95
rect 2097 51 2163 61
rect 2197 95 2251 111
rect 2197 61 2207 95
rect 2241 61 2251 95
rect 2197 17 2251 61
rect 2285 95 2351 129
rect 2473 129 2489 145
rect 2523 145 2677 163
rect 2523 129 2539 145
rect 2285 61 2301 95
rect 2335 61 2351 95
rect 2285 51 2351 61
rect 2385 95 2439 111
rect 2385 61 2395 95
rect 2429 61 2439 95
rect 2385 17 2439 61
rect 2473 95 2539 129
rect 2661 129 2677 145
rect 2711 145 2865 163
rect 2711 129 2727 145
rect 2473 61 2489 95
rect 2523 61 2539 95
rect 2473 51 2539 61
rect 2573 95 2627 111
rect 2573 61 2583 95
rect 2617 61 2627 95
rect 2573 17 2627 61
rect 2661 95 2727 129
rect 2849 129 2865 145
rect 2899 145 3053 163
rect 2899 129 2915 145
rect 2661 61 2677 95
rect 2711 61 2727 95
rect 2661 51 2727 61
rect 2761 95 2815 111
rect 2761 61 2771 95
rect 2805 61 2815 95
rect 2761 17 2815 61
rect 2849 95 2915 129
rect 3037 129 3053 145
rect 3087 129 3103 163
rect 2849 61 2865 95
rect 2899 61 2915 95
rect 2849 51 2915 61
rect 2949 95 3003 111
rect 2949 61 2961 95
rect 2995 61 3003 95
rect 2949 17 3003 61
rect 3037 95 3103 129
rect 3037 61 3053 95
rect 3087 61 3103 95
rect 3037 51 3103 61
rect 3137 163 3193 181
rect 3137 129 3149 163
rect 3183 129 3193 163
rect 3137 95 3193 129
rect 3137 61 3149 95
rect 3183 61 3193 95
rect 3137 17 3193 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3220 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
<< metal1 >>
rect 0 561 3220 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3220 561
rect 0 496 3220 527
rect 0 17 3220 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3220 17
rect 0 -48 3220 -17
<< labels >>
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 2053 221 2087 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 2881 221 2915 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 2513 221 2547 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4_8
<< properties >>
string FIXED_BBOX 0 0 3220 544
string GDS_END 405250
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 381744
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
