magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 53 21 907 203
rect 53 17 64 21
rect 30 -17 64 17
<< scnmos >>
rect 141 47 171 177
rect 235 47 265 177
rect 319 47 349 177
rect 413 47 443 177
rect 507 47 537 177
rect 601 47 631 177
rect 695 47 725 177
rect 799 47 829 177
<< scpmoshvt >>
rect 133 297 169 497
rect 227 297 263 497
rect 321 297 357 497
rect 415 297 451 497
rect 509 297 545 497
rect 603 297 639 497
rect 697 297 733 497
rect 791 297 827 497
<< ndiff >>
rect 79 97 141 177
rect 79 63 87 97
rect 121 63 141 97
rect 79 47 141 63
rect 171 161 235 177
rect 171 127 181 161
rect 215 127 235 161
rect 171 93 235 127
rect 171 59 181 93
rect 215 59 235 93
rect 171 47 235 59
rect 265 97 319 177
rect 265 63 275 97
rect 309 63 319 97
rect 265 47 319 63
rect 349 129 413 177
rect 349 95 369 129
rect 403 95 413 129
rect 349 47 413 95
rect 443 97 507 177
rect 443 63 463 97
rect 497 63 507 97
rect 443 47 507 63
rect 537 129 601 177
rect 537 95 557 129
rect 591 95 601 129
rect 537 47 601 95
rect 631 97 695 177
rect 631 63 651 97
rect 685 63 695 97
rect 631 47 695 63
rect 725 129 799 177
rect 725 95 745 129
rect 779 95 799 129
rect 725 47 799 95
rect 829 161 881 177
rect 829 127 839 161
rect 873 127 881 161
rect 829 93 881 127
rect 829 59 839 93
rect 873 59 881 93
rect 829 47 881 59
<< pdiff >>
rect 79 485 133 497
rect 79 451 87 485
rect 121 451 133 485
rect 79 417 133 451
rect 79 383 87 417
rect 121 383 133 417
rect 79 349 133 383
rect 79 315 87 349
rect 121 315 133 349
rect 79 297 133 315
rect 169 479 227 497
rect 169 445 181 479
rect 215 445 227 479
rect 169 411 227 445
rect 169 377 181 411
rect 215 377 227 411
rect 169 343 227 377
rect 169 309 181 343
rect 215 309 227 343
rect 169 297 227 309
rect 263 485 321 497
rect 263 451 275 485
rect 309 451 321 485
rect 263 417 321 451
rect 263 383 275 417
rect 309 383 321 417
rect 263 297 321 383
rect 357 463 415 497
rect 357 429 369 463
rect 403 429 415 463
rect 357 368 415 429
rect 357 334 369 368
rect 403 334 415 368
rect 357 297 415 334
rect 451 485 509 497
rect 451 451 463 485
rect 497 451 509 485
rect 451 417 509 451
rect 451 383 463 417
rect 497 383 509 417
rect 451 297 509 383
rect 545 463 603 497
rect 545 429 557 463
rect 591 429 603 463
rect 545 368 603 429
rect 545 334 557 368
rect 591 334 603 368
rect 545 297 603 334
rect 639 485 697 497
rect 639 451 651 485
rect 685 451 697 485
rect 639 417 697 451
rect 639 383 651 417
rect 685 383 697 417
rect 639 297 697 383
rect 733 463 791 497
rect 733 429 745 463
rect 779 429 791 463
rect 733 368 791 429
rect 733 334 745 368
rect 779 334 791 368
rect 733 297 791 334
rect 827 485 881 497
rect 827 451 839 485
rect 873 451 881 485
rect 827 417 881 451
rect 827 383 839 417
rect 873 383 881 417
rect 827 349 881 383
rect 827 315 839 349
rect 873 315 881 349
rect 827 297 881 315
<< ndiffc >>
rect 87 63 121 97
rect 181 127 215 161
rect 181 59 215 93
rect 275 63 309 97
rect 369 95 403 129
rect 463 63 497 97
rect 557 95 591 129
rect 651 63 685 97
rect 745 95 779 129
rect 839 127 873 161
rect 839 59 873 93
<< pdiffc >>
rect 87 451 121 485
rect 87 383 121 417
rect 87 315 121 349
rect 181 445 215 479
rect 181 377 215 411
rect 181 309 215 343
rect 275 451 309 485
rect 275 383 309 417
rect 369 429 403 463
rect 369 334 403 368
rect 463 451 497 485
rect 463 383 497 417
rect 557 429 591 463
rect 557 334 591 368
rect 651 451 685 485
rect 651 383 685 417
rect 745 429 779 463
rect 745 334 779 368
rect 839 451 873 485
rect 839 383 873 417
rect 839 315 873 349
<< poly >>
rect 133 497 169 523
rect 227 497 263 523
rect 321 497 357 523
rect 415 497 451 523
rect 509 497 545 523
rect 603 497 639 523
rect 697 497 733 523
rect 791 497 827 523
rect 133 282 169 297
rect 227 282 263 297
rect 321 282 357 297
rect 415 282 451 297
rect 509 282 545 297
rect 603 282 639 297
rect 697 282 733 297
rect 791 282 827 297
rect 131 259 171 282
rect 225 259 265 282
rect 65 249 265 259
rect 65 215 92 249
rect 126 215 197 249
rect 231 215 265 249
rect 65 205 265 215
rect 141 177 171 205
rect 235 177 265 205
rect 319 259 359 282
rect 413 259 453 282
rect 507 259 547 282
rect 601 259 641 282
rect 695 259 735 282
rect 789 259 829 282
rect 319 249 829 259
rect 319 215 335 249
rect 369 215 829 249
rect 319 205 829 215
rect 319 177 349 205
rect 413 177 443 205
rect 507 177 537 205
rect 601 177 631 205
rect 695 177 725 205
rect 799 177 829 205
rect 141 21 171 47
rect 235 21 265 47
rect 319 21 349 47
rect 413 21 443 47
rect 507 21 537 47
rect 601 21 631 47
rect 695 21 725 47
rect 799 21 829 47
<< polycont >>
rect 92 215 126 249
rect 197 215 231 249
rect 335 215 369 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 87 485 121 527
rect 87 417 121 451
rect 87 349 121 383
rect 87 297 121 315
rect 155 479 231 493
rect 155 445 181 479
rect 215 445 231 479
rect 155 411 231 445
rect 155 377 181 411
rect 215 377 231 411
rect 155 343 231 377
rect 275 485 323 527
rect 309 451 323 485
rect 275 417 323 451
rect 309 383 323 417
rect 275 367 323 383
rect 369 463 403 493
rect 369 368 403 429
rect 155 309 181 343
rect 215 331 231 343
rect 437 485 513 527
rect 437 451 463 485
rect 497 451 513 485
rect 437 417 513 451
rect 437 383 463 417
rect 497 383 513 417
rect 437 367 513 383
rect 557 463 591 493
rect 557 368 591 429
rect 215 309 325 331
rect 155 297 325 309
rect 56 249 253 263
rect 56 215 92 249
rect 126 215 197 249
rect 231 215 253 249
rect 291 249 325 297
rect 369 323 403 334
rect 625 485 701 527
rect 625 451 651 485
rect 685 451 701 485
rect 625 417 701 451
rect 625 383 651 417
rect 685 383 701 417
rect 625 367 701 383
rect 745 463 779 493
rect 745 368 779 429
rect 557 323 591 334
rect 745 323 779 334
rect 369 289 779 323
rect 813 485 889 527
rect 813 451 839 485
rect 873 451 889 485
rect 813 417 889 451
rect 813 383 839 417
rect 873 383 889 417
rect 813 349 889 383
rect 813 315 839 349
rect 873 315 889 349
rect 813 297 889 315
rect 291 215 335 249
rect 369 215 395 249
rect 291 181 325 215
rect 482 181 779 289
rect 155 161 325 181
rect 155 127 181 161
rect 215 147 325 161
rect 369 147 779 181
rect 215 127 231 147
rect 87 97 121 113
rect 87 17 121 63
rect 155 93 231 127
rect 369 129 403 147
rect 155 59 181 93
rect 215 59 231 93
rect 155 51 231 59
rect 275 97 309 113
rect 275 17 309 63
rect 557 129 591 147
rect 369 51 403 95
rect 437 97 513 113
rect 437 63 463 97
rect 497 63 513 97
rect 437 17 513 63
rect 745 129 779 147
rect 557 51 591 95
rect 625 97 701 113
rect 625 63 651 97
rect 685 63 701 97
rect 625 17 701 63
rect 745 51 779 95
rect 813 161 889 177
rect 813 127 839 161
rect 873 127 889 161
rect 813 93 889 127
rect 813 59 839 93
rect 873 59 889 93
rect 813 17 889 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 505 221 539 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 505 289 539 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 505 153 539 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional
flabel locali s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 188 221 222 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 78 221 112 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 buf_6
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 950836
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 943442
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
