magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1913 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 173 47 203 177
rect 267 47 297 177
rect 371 47 401 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 747 47 777 177
rect 935 47 965 177
rect 1029 47 1059 177
rect 1123 47 1153 177
rect 1227 47 1257 177
rect 1311 47 1341 177
rect 1405 47 1435 177
rect 1499 47 1529 177
rect 1593 47 1623 177
rect 1791 47 1821 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1125 297 1161 497
rect 1219 297 1255 497
rect 1313 297 1349 497
rect 1407 297 1443 497
rect 1501 297 1537 497
rect 1595 297 1631 497
rect 1793 297 1829 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 173 177
rect 109 129 129 163
rect 163 129 173 163
rect 109 95 173 129
rect 109 61 129 95
rect 163 61 173 95
rect 109 47 173 61
rect 203 95 267 177
rect 203 61 223 95
rect 257 61 267 95
rect 203 47 267 61
rect 297 163 371 177
rect 297 129 317 163
rect 351 129 371 163
rect 297 95 371 129
rect 297 61 317 95
rect 351 61 371 95
rect 297 47 371 61
rect 401 95 455 177
rect 401 61 411 95
rect 445 61 455 95
rect 401 47 455 61
rect 485 163 549 177
rect 485 129 505 163
rect 539 129 549 163
rect 485 95 549 129
rect 485 61 505 95
rect 539 61 549 95
rect 485 47 549 61
rect 579 95 643 177
rect 579 61 599 95
rect 633 61 643 95
rect 579 47 643 61
rect 673 163 747 177
rect 673 129 693 163
rect 727 129 747 163
rect 673 95 747 129
rect 673 61 693 95
rect 727 61 747 95
rect 673 47 747 61
rect 777 95 935 177
rect 777 61 787 95
rect 821 61 891 95
rect 925 61 935 95
rect 777 47 935 61
rect 965 163 1029 177
rect 965 129 985 163
rect 1019 129 1029 163
rect 965 95 1029 129
rect 965 61 985 95
rect 1019 61 1029 95
rect 965 47 1029 61
rect 1059 95 1123 177
rect 1059 61 1079 95
rect 1113 61 1123 95
rect 1059 47 1123 61
rect 1153 163 1227 177
rect 1153 129 1173 163
rect 1207 129 1227 163
rect 1153 95 1227 129
rect 1153 61 1173 95
rect 1207 61 1227 95
rect 1153 47 1227 61
rect 1257 95 1311 177
rect 1257 61 1267 95
rect 1301 61 1311 95
rect 1257 47 1311 61
rect 1341 163 1405 177
rect 1341 129 1361 163
rect 1395 129 1405 163
rect 1341 95 1405 129
rect 1341 61 1361 95
rect 1395 61 1405 95
rect 1341 47 1405 61
rect 1435 95 1499 177
rect 1435 61 1455 95
rect 1489 61 1499 95
rect 1435 47 1499 61
rect 1529 163 1593 177
rect 1529 129 1549 163
rect 1583 129 1593 163
rect 1529 95 1593 129
rect 1529 61 1549 95
rect 1583 61 1593 95
rect 1529 47 1593 61
rect 1623 95 1685 177
rect 1623 61 1643 95
rect 1677 61 1685 95
rect 1623 47 1685 61
rect 1739 163 1791 177
rect 1739 129 1747 163
rect 1781 129 1791 163
rect 1739 95 1791 129
rect 1739 61 1747 95
rect 1781 61 1791 95
rect 1739 47 1791 61
rect 1821 163 1887 177
rect 1821 129 1841 163
rect 1875 129 1887 163
rect 1821 95 1887 129
rect 1821 61 1841 95
rect 1875 61 1887 95
rect 1821 47 1887 61
<< pdiff >>
rect 27 479 81 497
rect 27 445 35 479
rect 69 445 81 479
rect 27 411 81 445
rect 27 377 35 411
rect 69 377 81 411
rect 27 343 81 377
rect 27 309 35 343
rect 69 309 81 343
rect 27 297 81 309
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 297 175 375
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 409 269 443
rect 211 375 223 409
rect 257 375 269 409
rect 211 341 269 375
rect 211 307 223 341
rect 257 307 269 341
rect 211 297 269 307
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 409 363 443
rect 305 375 317 409
rect 351 375 363 409
rect 305 297 363 375
rect 399 477 457 497
rect 399 443 411 477
rect 445 443 457 477
rect 399 409 457 443
rect 399 375 411 409
rect 445 375 457 409
rect 399 341 457 375
rect 399 307 411 341
rect 445 307 457 341
rect 399 297 457 307
rect 493 409 551 497
rect 493 375 505 409
rect 539 375 551 409
rect 493 341 551 375
rect 493 307 505 341
rect 539 307 551 341
rect 493 297 551 307
rect 587 477 645 497
rect 587 443 599 477
rect 633 443 645 477
rect 587 409 645 443
rect 587 375 599 409
rect 633 375 645 409
rect 587 297 645 375
rect 681 409 739 497
rect 681 375 693 409
rect 727 375 739 409
rect 681 341 739 375
rect 681 307 693 341
rect 727 307 739 341
rect 681 297 739 307
rect 775 477 829 497
rect 775 443 787 477
rect 821 443 829 477
rect 775 409 829 443
rect 775 375 787 409
rect 821 375 829 409
rect 775 297 829 375
rect 883 477 937 497
rect 883 443 891 477
rect 925 443 937 477
rect 883 409 937 443
rect 883 375 891 409
rect 925 375 937 409
rect 883 297 937 375
rect 973 409 1031 497
rect 973 375 985 409
rect 1019 375 1031 409
rect 973 341 1031 375
rect 973 307 985 341
rect 1019 307 1031 341
rect 973 297 1031 307
rect 1067 477 1125 497
rect 1067 443 1079 477
rect 1113 443 1125 477
rect 1067 409 1125 443
rect 1067 375 1079 409
rect 1113 375 1125 409
rect 1067 297 1125 375
rect 1161 409 1219 497
rect 1161 375 1173 409
rect 1207 375 1219 409
rect 1161 341 1219 375
rect 1161 307 1173 341
rect 1207 307 1219 341
rect 1161 297 1219 307
rect 1255 477 1313 497
rect 1255 443 1267 477
rect 1301 443 1313 477
rect 1255 409 1313 443
rect 1255 375 1267 409
rect 1301 375 1313 409
rect 1255 341 1313 375
rect 1255 307 1267 341
rect 1301 307 1313 341
rect 1255 297 1313 307
rect 1349 409 1407 497
rect 1349 375 1361 409
rect 1395 375 1407 409
rect 1349 341 1407 375
rect 1349 307 1361 341
rect 1395 307 1407 341
rect 1349 297 1407 307
rect 1443 477 1501 497
rect 1443 443 1455 477
rect 1489 443 1501 477
rect 1443 409 1501 443
rect 1443 375 1455 409
rect 1489 375 1501 409
rect 1443 297 1501 375
rect 1537 409 1595 497
rect 1537 375 1549 409
rect 1583 375 1595 409
rect 1537 341 1595 375
rect 1537 307 1549 341
rect 1583 307 1595 341
rect 1537 297 1595 307
rect 1631 477 1685 497
rect 1631 443 1643 477
rect 1677 443 1685 477
rect 1631 409 1685 443
rect 1631 375 1643 409
rect 1677 375 1685 409
rect 1631 297 1685 375
rect 1739 479 1793 497
rect 1739 445 1747 479
rect 1781 445 1793 479
rect 1739 411 1793 445
rect 1739 377 1747 411
rect 1781 377 1793 411
rect 1739 343 1793 377
rect 1739 309 1747 343
rect 1781 309 1793 343
rect 1739 297 1793 309
rect 1829 479 1887 497
rect 1829 445 1841 479
rect 1875 445 1887 479
rect 1829 411 1887 445
rect 1829 377 1841 411
rect 1875 377 1887 411
rect 1829 343 1887 377
rect 1829 309 1841 343
rect 1875 309 1887 343
rect 1829 297 1887 309
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 129 129 163 163
rect 129 61 163 95
rect 223 61 257 95
rect 317 129 351 163
rect 317 61 351 95
rect 411 61 445 95
rect 505 129 539 163
rect 505 61 539 95
rect 599 61 633 95
rect 693 129 727 163
rect 693 61 727 95
rect 787 61 821 95
rect 891 61 925 95
rect 985 129 1019 163
rect 985 61 1019 95
rect 1079 61 1113 95
rect 1173 129 1207 163
rect 1173 61 1207 95
rect 1267 61 1301 95
rect 1361 129 1395 163
rect 1361 61 1395 95
rect 1455 61 1489 95
rect 1549 129 1583 163
rect 1549 61 1583 95
rect 1643 61 1677 95
rect 1747 129 1781 163
rect 1747 61 1781 95
rect 1841 129 1875 163
rect 1841 61 1875 95
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 129 443 163 477
rect 129 375 163 409
rect 223 443 257 477
rect 223 375 257 409
rect 223 307 257 341
rect 317 443 351 477
rect 317 375 351 409
rect 411 443 445 477
rect 411 375 445 409
rect 411 307 445 341
rect 505 375 539 409
rect 505 307 539 341
rect 599 443 633 477
rect 599 375 633 409
rect 693 375 727 409
rect 693 307 727 341
rect 787 443 821 477
rect 787 375 821 409
rect 891 443 925 477
rect 891 375 925 409
rect 985 375 1019 409
rect 985 307 1019 341
rect 1079 443 1113 477
rect 1079 375 1113 409
rect 1173 375 1207 409
rect 1173 307 1207 341
rect 1267 443 1301 477
rect 1267 375 1301 409
rect 1267 307 1301 341
rect 1361 375 1395 409
rect 1361 307 1395 341
rect 1455 443 1489 477
rect 1455 375 1489 409
rect 1549 375 1583 409
rect 1549 307 1583 341
rect 1643 443 1677 477
rect 1643 375 1677 409
rect 1747 445 1781 479
rect 1747 377 1781 411
rect 1747 309 1781 343
rect 1841 445 1875 479
rect 1841 377 1875 411
rect 1841 309 1875 343
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1125 497 1161 523
rect 1219 497 1255 523
rect 1313 497 1349 523
rect 1407 497 1443 523
rect 1501 497 1537 523
rect 1595 497 1631 523
rect 1793 497 1829 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1125 282 1161 297
rect 1219 282 1255 297
rect 1313 282 1349 297
rect 1407 282 1443 297
rect 1501 282 1537 297
rect 1595 282 1631 297
rect 1793 282 1829 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 79 249 401 265
rect 79 215 95 249
rect 129 215 173 249
rect 207 215 251 249
rect 285 215 329 249
rect 363 215 401 249
rect 79 199 401 215
rect 79 177 109 199
rect 173 177 203 199
rect 267 177 297 199
rect 371 177 401 199
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 455 249 777 265
rect 455 215 471 249
rect 505 215 549 249
rect 583 215 627 249
rect 661 215 705 249
rect 739 215 777 249
rect 455 199 777 215
rect 455 177 485 199
rect 549 177 579 199
rect 643 177 673 199
rect 747 177 777 199
rect 935 265 975 282
rect 1029 265 1069 282
rect 1123 265 1163 282
rect 1217 265 1257 282
rect 935 249 1257 265
rect 935 215 951 249
rect 985 215 1029 249
rect 1063 215 1107 249
rect 1141 215 1185 249
rect 1219 215 1257 249
rect 935 199 1257 215
rect 935 177 965 199
rect 1029 177 1059 199
rect 1123 177 1153 199
rect 1227 177 1257 199
rect 1311 265 1351 282
rect 1405 265 1445 282
rect 1499 265 1539 282
rect 1593 265 1633 282
rect 1791 265 1831 282
rect 1311 249 1704 265
rect 1311 215 1508 249
rect 1542 215 1586 249
rect 1620 215 1654 249
rect 1688 215 1704 249
rect 1311 199 1704 215
rect 1791 249 1882 265
rect 1791 215 1832 249
rect 1866 215 1882 249
rect 1791 199 1882 215
rect 1311 177 1341 199
rect 1405 177 1435 199
rect 1499 177 1529 199
rect 1593 177 1623 199
rect 1791 177 1821 199
rect 79 21 109 47
rect 173 21 203 47
rect 267 21 297 47
rect 371 21 401 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 747 21 777 47
rect 935 21 965 47
rect 1029 21 1059 47
rect 1123 21 1153 47
rect 1227 21 1257 47
rect 1311 21 1341 47
rect 1405 21 1435 47
rect 1499 21 1529 47
rect 1593 21 1623 47
rect 1791 21 1821 47
<< polycont >>
rect 95 215 129 249
rect 173 215 207 249
rect 251 215 285 249
rect 329 215 363 249
rect 471 215 505 249
rect 549 215 583 249
rect 627 215 661 249
rect 705 215 739 249
rect 951 215 985 249
rect 1029 215 1063 249
rect 1107 215 1141 249
rect 1185 215 1219 249
rect 1508 215 1542 249
rect 1586 215 1620 249
rect 1654 215 1688 249
rect 1832 215 1866 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 19 479 85 493
rect 19 445 35 479
rect 69 445 85 479
rect 19 411 85 445
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 129 477 171 527
rect 163 443 171 477
rect 129 409 171 443
rect 163 375 171 409
rect 129 359 171 375
rect 215 477 265 493
rect 215 443 223 477
rect 257 443 265 477
rect 215 409 265 443
rect 215 375 223 409
rect 257 375 265 409
rect 19 309 35 343
rect 69 325 85 343
rect 215 341 265 375
rect 309 477 359 527
rect 309 443 317 477
rect 351 443 359 477
rect 309 409 359 443
rect 309 375 317 409
rect 351 375 359 409
rect 309 359 359 375
rect 403 477 829 493
rect 403 443 411 477
rect 445 459 599 477
rect 445 443 453 459
rect 403 409 453 443
rect 591 443 599 459
rect 633 459 787 477
rect 633 443 641 459
rect 403 375 411 409
rect 445 375 453 409
rect 215 325 223 341
rect 69 309 223 325
rect 19 307 223 309
rect 257 325 265 341
rect 403 341 453 375
rect 403 325 411 341
rect 257 307 411 325
rect 445 307 453 341
rect 19 291 453 307
rect 497 409 547 425
rect 497 375 505 409
rect 539 375 547 409
rect 497 341 547 375
rect 591 409 641 443
rect 779 443 787 459
rect 821 443 829 477
rect 591 375 599 409
rect 633 375 641 409
rect 591 359 641 375
rect 685 409 735 425
rect 685 375 693 409
rect 727 375 735 409
rect 497 307 505 341
rect 539 325 547 341
rect 685 341 735 375
rect 779 409 829 443
rect 779 375 787 409
rect 821 375 829 409
rect 779 359 829 375
rect 883 477 1685 493
rect 883 443 891 477
rect 925 459 1079 477
rect 925 443 933 459
rect 883 409 933 443
rect 1071 443 1079 459
rect 1113 459 1267 477
rect 1113 443 1121 459
rect 883 375 891 409
rect 925 375 933 409
rect 883 359 933 375
rect 977 409 1027 425
rect 977 375 985 409
rect 1019 375 1027 409
rect 685 325 693 341
rect 539 307 693 325
rect 727 325 735 341
rect 977 341 1027 375
rect 1071 409 1121 443
rect 1259 443 1267 459
rect 1301 459 1455 477
rect 1301 443 1309 459
rect 1071 375 1079 409
rect 1113 375 1121 409
rect 1071 359 1121 375
rect 1165 409 1215 425
rect 1165 375 1173 409
rect 1207 375 1215 409
rect 977 325 985 341
rect 727 307 985 325
rect 1019 325 1027 341
rect 1165 341 1215 375
rect 1165 325 1173 341
rect 1019 307 1173 325
rect 1207 307 1215 341
rect 497 291 1215 307
rect 1259 409 1309 443
rect 1447 443 1455 459
rect 1489 459 1643 477
rect 1489 443 1497 459
rect 1259 375 1267 409
rect 1301 375 1309 409
rect 1259 341 1309 375
rect 1259 307 1267 341
rect 1301 307 1309 341
rect 1259 291 1309 307
rect 1353 409 1403 425
rect 1353 375 1361 409
rect 1395 375 1403 409
rect 1353 341 1403 375
rect 1447 409 1497 443
rect 1635 443 1643 459
rect 1677 443 1685 477
rect 1447 375 1455 409
rect 1489 375 1497 409
rect 1447 359 1497 375
rect 1541 409 1591 425
rect 1541 375 1549 409
rect 1583 375 1591 409
rect 1353 307 1361 341
rect 1395 325 1403 341
rect 1541 341 1591 375
rect 1635 409 1685 443
rect 1635 375 1643 409
rect 1677 375 1685 409
rect 1635 359 1685 375
rect 1730 479 1797 493
rect 1730 445 1747 479
rect 1781 445 1797 479
rect 1730 411 1797 445
rect 1730 377 1747 411
rect 1781 377 1797 411
rect 1541 325 1549 341
rect 1395 307 1549 325
rect 1583 307 1591 341
rect 1730 343 1797 377
rect 1730 325 1747 343
rect 1353 291 1591 307
rect 1654 309 1747 325
rect 1781 309 1797 343
rect 1654 291 1797 309
rect 1841 479 1887 527
rect 1875 445 1887 479
rect 1841 411 1887 445
rect 1875 377 1887 411
rect 1841 343 1887 377
rect 1875 309 1887 343
rect 1841 291 1887 309
rect 79 249 401 257
rect 79 215 95 249
rect 129 215 173 249
rect 207 215 251 249
rect 285 215 329 249
rect 363 215 401 249
rect 455 249 830 257
rect 455 215 471 249
rect 505 215 549 249
rect 583 215 627 249
rect 661 215 705 249
rect 739 215 830 249
rect 877 249 1257 257
rect 877 215 951 249
rect 985 215 1029 249
rect 1063 215 1107 249
rect 1141 215 1185 249
rect 1219 215 1257 249
rect 1353 181 1450 291
rect 1654 257 1688 291
rect 1484 249 1688 257
rect 1484 215 1508 249
rect 1542 215 1586 249
rect 1620 215 1654 249
rect 1771 249 1910 257
rect 1771 215 1832 249
rect 1866 215 1910 249
rect 1654 181 1688 215
rect 35 163 69 179
rect 35 95 69 129
rect 35 17 69 61
rect 103 163 1599 181
rect 103 129 129 163
rect 163 145 317 163
rect 163 129 179 145
rect 103 95 179 129
rect 291 129 317 145
rect 351 145 505 163
rect 351 129 367 145
rect 103 61 129 95
rect 163 61 179 95
rect 103 51 179 61
rect 223 95 257 111
rect 223 17 257 61
rect 291 95 367 129
rect 479 129 505 145
rect 539 145 693 163
rect 539 129 555 145
rect 291 61 317 95
rect 351 61 367 95
rect 291 51 367 61
rect 411 95 445 111
rect 411 17 445 61
rect 479 95 555 129
rect 667 129 693 145
rect 727 145 985 163
rect 727 129 743 145
rect 479 61 505 95
rect 539 61 555 95
rect 479 51 555 61
rect 599 95 633 111
rect 599 17 633 61
rect 667 95 743 129
rect 959 129 985 145
rect 1019 145 1173 163
rect 1019 129 1035 145
rect 667 61 693 95
rect 727 61 743 95
rect 667 51 743 61
rect 787 95 925 111
rect 821 61 891 95
rect 787 17 925 61
rect 959 95 1035 129
rect 1147 129 1173 145
rect 1207 145 1361 163
rect 1207 129 1223 145
rect 959 61 985 95
rect 1019 61 1035 95
rect 959 51 1035 61
rect 1079 95 1113 111
rect 1079 17 1113 61
rect 1147 95 1223 129
rect 1335 129 1361 145
rect 1395 145 1549 163
rect 1395 129 1411 145
rect 1147 61 1173 95
rect 1207 61 1223 95
rect 1147 51 1223 61
rect 1267 95 1301 111
rect 1267 17 1301 61
rect 1335 95 1411 129
rect 1523 129 1549 145
rect 1583 129 1599 163
rect 1654 163 1797 181
rect 1654 147 1747 163
rect 1335 61 1361 95
rect 1395 61 1411 95
rect 1335 51 1411 61
rect 1455 95 1489 111
rect 1455 17 1489 61
rect 1523 95 1599 129
rect 1722 129 1747 147
rect 1781 129 1797 163
rect 1523 61 1549 95
rect 1583 61 1599 95
rect 1523 51 1599 61
rect 1643 95 1677 111
rect 1643 17 1677 61
rect 1722 95 1797 129
rect 1722 61 1747 95
rect 1781 61 1797 95
rect 1722 51 1797 61
rect 1841 163 1887 181
rect 1875 129 1887 163
rect 1841 95 1887 129
rect 1875 61 1887 95
rect 1841 17 1887 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 455 215 830 257 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 79 215 401 257 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 1856 221 1890 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 1039 221 1075 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 1356 357 1390 391 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4b_4
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_END 1819346
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1805020
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
