magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 5 21 295 203
rect 28 -17 62 21
<< scnmos >>
rect 93 47 123 177
rect 177 47 207 177
<< scpmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
<< ndiff >>
rect 31 161 93 177
rect 31 127 39 161
rect 73 127 93 161
rect 31 93 93 127
rect 31 59 39 93
rect 73 59 93 93
rect 31 47 93 59
rect 123 47 177 177
rect 207 161 269 177
rect 207 127 227 161
rect 261 127 269 161
rect 207 93 269 127
rect 207 59 227 93
rect 261 59 269 93
rect 207 47 269 59
<< pdiff >>
rect 31 485 85 497
rect 31 451 39 485
rect 73 451 85 485
rect 31 417 85 451
rect 31 383 39 417
rect 73 383 85 417
rect 31 349 85 383
rect 31 315 39 349
rect 73 315 85 349
rect 31 297 85 315
rect 121 485 179 497
rect 121 451 133 485
rect 167 451 179 485
rect 121 417 179 451
rect 121 383 133 417
rect 167 383 179 417
rect 121 349 179 383
rect 121 315 133 349
rect 167 315 179 349
rect 121 297 179 315
rect 215 485 269 497
rect 215 451 227 485
rect 261 451 269 485
rect 215 417 269 451
rect 215 383 227 417
rect 261 383 269 417
rect 215 349 269 383
rect 215 315 227 349
rect 261 315 269 349
rect 215 297 269 315
<< ndiffc >>
rect 39 127 73 161
rect 39 59 73 93
rect 227 127 261 161
rect 227 59 261 93
<< pdiffc >>
rect 39 451 73 485
rect 39 383 73 417
rect 39 315 73 349
rect 133 451 167 485
rect 133 383 167 417
rect 133 315 167 349
rect 227 451 261 485
rect 227 383 261 417
rect 227 315 261 349
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 85 282 121 297
rect 179 282 215 297
rect 83 265 123 282
rect 21 249 123 265
rect 21 215 36 249
rect 70 215 123 249
rect 21 199 123 215
rect 93 177 123 199
rect 177 265 217 282
rect 177 249 275 265
rect 177 215 224 249
rect 258 215 275 249
rect 177 199 275 215
rect 177 177 207 199
rect 93 21 123 47
rect 177 21 207 47
<< polycont >>
rect 36 215 70 249
rect 224 215 258 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 17 485 73 527
rect 17 451 39 485
rect 17 417 73 451
rect 17 383 39 417
rect 17 349 73 383
rect 17 315 39 349
rect 17 299 73 315
rect 107 485 183 493
rect 107 451 133 485
rect 167 451 183 485
rect 107 417 183 451
rect 107 383 133 417
rect 167 383 183 417
rect 107 349 183 383
rect 107 315 133 349
rect 167 315 183 349
rect 107 297 183 315
rect 227 485 279 527
rect 261 451 279 485
rect 227 417 279 451
rect 261 383 279 417
rect 227 349 279 383
rect 261 315 279 349
rect 227 299 279 315
rect 19 249 86 265
rect 19 215 36 249
rect 70 215 86 249
rect 19 211 86 215
rect 130 177 164 297
rect 198 249 275 265
rect 198 215 224 249
rect 258 215 275 249
rect 17 161 79 177
rect 17 127 39 161
rect 73 127 79 161
rect 17 93 79 127
rect 17 59 39 93
rect 73 59 79 93
rect 17 17 79 59
rect 130 161 279 177
rect 130 127 227 161
rect 261 127 279 161
rect 130 93 279 127
rect 130 59 227 93
rect 261 59 279 93
rect 130 51 279 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel locali s 130 296 164 330 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 130 364 164 398 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 212 141 246 175 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 28 221 62 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 198 215 275 265 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel nwell s 28 527 62 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 28 -17 62 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 28 -17 62 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 28 527 62 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2_1
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_END 1480002
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1475886
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
