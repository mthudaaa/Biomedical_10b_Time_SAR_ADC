magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 1 21 2107 203
rect 30 -17 64 21
<< scnmos >>
rect 93 47 123 177
rect 187 47 217 177
rect 281 47 311 177
rect 375 47 405 177
rect 573 47 603 177
rect 667 47 697 177
rect 761 47 791 177
rect 845 47 875 177
rect 939 47 969 177
rect 1033 47 1063 177
rect 1137 47 1167 177
rect 1231 47 1261 177
rect 1341 47 1371 177
rect 1425 47 1455 177
rect 1519 47 1549 177
rect 1613 47 1643 177
rect 1717 47 1747 177
rect 1801 47 1831 177
rect 1895 47 1925 177
rect 1989 47 2019 177
<< scpmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 565 297 601 497
rect 659 297 695 497
rect 753 297 789 497
rect 847 297 883 497
rect 941 297 977 497
rect 1035 297 1071 497
rect 1129 297 1165 497
rect 1223 297 1259 497
rect 1333 297 1369 497
rect 1427 297 1463 497
rect 1521 297 1557 497
rect 1615 297 1651 497
rect 1709 297 1745 497
rect 1803 297 1839 497
rect 1897 297 1933 497
rect 1991 297 2027 497
<< ndiff >>
rect 27 163 93 177
rect 27 129 39 163
rect 73 129 93 163
rect 27 95 93 129
rect 27 61 39 95
rect 73 61 93 95
rect 27 47 93 61
rect 123 163 187 177
rect 123 129 133 163
rect 167 129 187 163
rect 123 47 187 129
rect 217 95 281 177
rect 217 61 227 95
rect 261 61 281 95
rect 217 47 281 61
rect 311 163 375 177
rect 311 129 321 163
rect 355 129 375 163
rect 311 47 375 129
rect 405 95 457 177
rect 405 61 415 95
rect 449 61 457 95
rect 405 47 457 61
rect 511 163 573 177
rect 511 129 519 163
rect 553 129 573 163
rect 511 47 573 129
rect 603 95 667 177
rect 603 61 613 95
rect 647 61 667 95
rect 603 47 667 61
rect 697 163 761 177
rect 697 129 707 163
rect 741 129 761 163
rect 697 47 761 129
rect 791 95 845 177
rect 791 61 801 95
rect 835 61 845 95
rect 791 47 845 61
rect 875 163 939 177
rect 875 129 895 163
rect 929 129 939 163
rect 875 47 939 129
rect 969 95 1033 177
rect 969 61 989 95
rect 1023 61 1033 95
rect 969 47 1033 61
rect 1063 163 1137 177
rect 1063 129 1083 163
rect 1117 129 1137 163
rect 1063 47 1137 129
rect 1167 95 1231 177
rect 1167 61 1177 95
rect 1211 61 1231 95
rect 1167 47 1231 61
rect 1261 163 1341 177
rect 1261 129 1287 163
rect 1321 129 1341 163
rect 1261 95 1341 129
rect 1261 61 1287 95
rect 1321 61 1341 95
rect 1261 47 1341 61
rect 1371 95 1425 177
rect 1371 61 1381 95
rect 1415 61 1425 95
rect 1371 47 1425 61
rect 1455 163 1519 177
rect 1455 129 1475 163
rect 1509 129 1519 163
rect 1455 95 1519 129
rect 1455 61 1475 95
rect 1509 61 1519 95
rect 1455 47 1519 61
rect 1549 95 1613 177
rect 1549 61 1569 95
rect 1603 61 1613 95
rect 1549 47 1613 61
rect 1643 163 1717 177
rect 1643 129 1663 163
rect 1697 129 1717 163
rect 1643 95 1717 129
rect 1643 61 1663 95
rect 1697 61 1717 95
rect 1643 47 1717 61
rect 1747 95 1801 177
rect 1747 61 1757 95
rect 1791 61 1801 95
rect 1747 47 1801 61
rect 1831 163 1895 177
rect 1831 129 1851 163
rect 1885 129 1895 163
rect 1831 95 1895 129
rect 1831 61 1851 95
rect 1885 61 1895 95
rect 1831 47 1895 61
rect 1925 95 1989 177
rect 1925 61 1945 95
rect 1979 61 1989 95
rect 1925 47 1989 61
rect 2019 163 2081 177
rect 2019 129 2039 163
rect 2073 129 2081 163
rect 2019 95 2081 129
rect 2019 61 2039 95
rect 2073 61 2081 95
rect 2019 47 2081 61
<< pdiff >>
rect 27 483 85 497
rect 27 449 39 483
rect 73 449 85 483
rect 27 415 85 449
rect 27 381 39 415
rect 73 381 85 415
rect 27 347 85 381
rect 27 313 39 347
rect 73 313 85 347
rect 27 297 85 313
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 341 179 375
rect 121 307 133 341
rect 167 307 179 341
rect 121 297 179 307
rect 215 483 273 497
rect 215 449 227 483
rect 261 449 273 483
rect 215 415 273 449
rect 215 381 227 415
rect 261 381 273 415
rect 215 297 273 381
rect 309 477 367 497
rect 309 443 321 477
rect 355 443 367 477
rect 309 409 367 443
rect 309 375 321 409
rect 355 375 367 409
rect 309 341 367 375
rect 309 307 321 341
rect 355 307 367 341
rect 309 297 367 307
rect 403 477 565 497
rect 403 443 415 477
rect 449 443 519 477
rect 553 443 565 477
rect 403 297 565 443
rect 601 477 659 497
rect 601 443 613 477
rect 647 443 659 477
rect 601 409 659 443
rect 601 375 613 409
rect 647 375 659 409
rect 601 297 659 375
rect 695 477 753 497
rect 695 443 707 477
rect 741 443 753 477
rect 695 297 753 443
rect 789 477 847 497
rect 789 443 801 477
rect 835 443 847 477
rect 789 409 847 443
rect 789 375 801 409
rect 835 375 847 409
rect 789 297 847 375
rect 883 401 941 497
rect 883 367 895 401
rect 929 367 941 401
rect 883 297 941 367
rect 977 487 1035 497
rect 977 453 989 487
rect 1023 453 1035 487
rect 977 297 1035 453
rect 1071 401 1129 497
rect 1071 367 1083 401
rect 1117 367 1129 401
rect 1071 297 1129 367
rect 1165 487 1223 497
rect 1165 453 1177 487
rect 1211 453 1223 487
rect 1165 297 1223 453
rect 1259 487 1333 497
rect 1259 453 1279 487
rect 1313 453 1333 487
rect 1259 297 1333 453
rect 1369 487 1427 497
rect 1369 453 1381 487
rect 1415 453 1427 487
rect 1369 297 1427 453
rect 1463 401 1521 497
rect 1463 367 1475 401
rect 1509 367 1521 401
rect 1463 297 1521 367
rect 1557 487 1615 497
rect 1557 453 1569 487
rect 1603 453 1615 487
rect 1557 297 1615 453
rect 1651 401 1709 497
rect 1651 367 1663 401
rect 1697 367 1709 401
rect 1651 297 1709 367
rect 1745 477 1803 497
rect 1745 443 1757 477
rect 1791 443 1803 477
rect 1745 409 1803 443
rect 1745 375 1757 409
rect 1791 375 1803 409
rect 1745 297 1803 375
rect 1839 477 1897 497
rect 1839 443 1851 477
rect 1885 443 1897 477
rect 1839 297 1897 443
rect 1933 477 1991 497
rect 1933 443 1945 477
rect 1979 443 1991 477
rect 1933 409 1991 443
rect 1933 375 1945 409
rect 1979 375 1991 409
rect 1933 341 1991 375
rect 1933 307 1945 341
rect 1979 307 1991 341
rect 1933 297 1991 307
rect 2027 477 2088 497
rect 2027 443 2039 477
rect 2073 443 2088 477
rect 2027 409 2088 443
rect 2027 375 2039 409
rect 2073 375 2088 409
rect 2027 341 2088 375
rect 2027 307 2039 341
rect 2073 307 2088 341
rect 2027 297 2088 307
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 227 61 261 95
rect 321 129 355 163
rect 415 61 449 95
rect 519 129 553 163
rect 613 61 647 95
rect 707 129 741 163
rect 801 61 835 95
rect 895 129 929 163
rect 989 61 1023 95
rect 1083 129 1117 163
rect 1177 61 1211 95
rect 1287 129 1321 163
rect 1287 61 1321 95
rect 1381 61 1415 95
rect 1475 129 1509 163
rect 1475 61 1509 95
rect 1569 61 1603 95
rect 1663 129 1697 163
rect 1663 61 1697 95
rect 1757 61 1791 95
rect 1851 129 1885 163
rect 1851 61 1885 95
rect 1945 61 1979 95
rect 2039 129 2073 163
rect 2039 61 2073 95
<< pdiffc >>
rect 39 449 73 483
rect 39 381 73 415
rect 39 313 73 347
rect 133 443 167 477
rect 133 375 167 409
rect 133 307 167 341
rect 227 449 261 483
rect 227 381 261 415
rect 321 443 355 477
rect 321 375 355 409
rect 321 307 355 341
rect 415 443 449 477
rect 519 443 553 477
rect 613 443 647 477
rect 613 375 647 409
rect 707 443 741 477
rect 801 443 835 477
rect 801 375 835 409
rect 895 367 929 401
rect 989 453 1023 487
rect 1083 367 1117 401
rect 1177 453 1211 487
rect 1279 453 1313 487
rect 1381 453 1415 487
rect 1475 367 1509 401
rect 1569 453 1603 487
rect 1663 367 1697 401
rect 1757 443 1791 477
rect 1757 375 1791 409
rect 1851 443 1885 477
rect 1945 443 1979 477
rect 1945 375 1979 409
rect 1945 307 1979 341
rect 2039 443 2073 477
rect 2039 375 2073 409
rect 2039 307 2073 341
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 565 497 601 523
rect 659 497 695 523
rect 753 497 789 523
rect 847 497 883 523
rect 941 497 977 523
rect 1035 497 1071 523
rect 1129 497 1165 523
rect 1223 497 1259 523
rect 1333 497 1369 523
rect 1427 497 1463 523
rect 1521 497 1557 523
rect 1615 497 1651 523
rect 1709 497 1745 523
rect 1803 497 1839 523
rect 1897 497 1933 523
rect 1991 497 2027 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 565 282 601 297
rect 659 282 695 297
rect 753 282 789 297
rect 847 282 883 297
rect 941 282 977 297
rect 1035 282 1071 297
rect 1129 282 1165 297
rect 1223 282 1259 297
rect 1333 282 1369 297
rect 1427 282 1463 297
rect 1521 282 1557 297
rect 1615 282 1651 297
rect 1709 282 1745 297
rect 1803 282 1839 297
rect 1897 282 1933 297
rect 1991 282 2027 297
rect 83 265 123 282
rect 177 265 217 282
rect 271 265 311 282
rect 365 265 405 282
rect 563 265 603 282
rect 657 265 697 282
rect 751 265 791 282
rect 65 249 405 265
rect 65 215 81 249
rect 115 215 159 249
rect 193 215 237 249
rect 271 215 315 249
rect 349 215 405 249
rect 65 199 405 215
rect 554 249 791 265
rect 554 215 570 249
rect 604 215 648 249
rect 682 215 726 249
rect 760 215 791 249
rect 554 199 791 215
rect 93 177 123 199
rect 187 177 217 199
rect 281 177 311 199
rect 375 177 405 199
rect 573 177 603 199
rect 667 177 697 199
rect 761 177 791 199
rect 845 265 885 282
rect 939 265 979 282
rect 1033 265 1073 282
rect 1127 265 1167 282
rect 1221 265 1261 282
rect 1331 265 1371 282
rect 1425 265 1465 282
rect 1519 265 1559 282
rect 1613 265 1653 282
rect 1707 265 1747 282
rect 845 249 1167 265
rect 845 215 1035 249
rect 1069 215 1113 249
rect 1147 215 1167 249
rect 845 199 1167 215
rect 1209 249 1273 265
rect 1209 215 1219 249
rect 1253 215 1273 249
rect 1209 199 1273 215
rect 1319 249 1383 265
rect 1319 215 1329 249
rect 1363 215 1383 249
rect 1319 199 1383 215
rect 1425 249 1747 265
rect 1425 215 1519 249
rect 1553 215 1590 249
rect 1624 215 1675 249
rect 1709 215 1747 249
rect 1425 199 1747 215
rect 845 177 875 199
rect 939 177 969 199
rect 1033 177 1063 199
rect 1137 177 1167 199
rect 1231 177 1261 199
rect 1341 177 1371 199
rect 1425 177 1455 199
rect 1519 177 1549 199
rect 1613 177 1643 199
rect 1717 177 1747 199
rect 1801 265 1841 282
rect 1895 265 1935 282
rect 1989 265 2029 282
rect 1801 249 2038 265
rect 1801 215 1817 249
rect 1851 215 1895 249
rect 1929 215 1973 249
rect 2007 215 2038 249
rect 1801 199 2038 215
rect 1801 177 1831 199
rect 1895 177 1925 199
rect 1989 177 2019 199
rect 93 21 123 47
rect 187 21 217 47
rect 281 21 311 47
rect 375 21 405 47
rect 573 21 603 47
rect 667 21 697 47
rect 761 21 791 47
rect 845 21 875 47
rect 939 21 969 47
rect 1033 21 1063 47
rect 1137 21 1167 47
rect 1231 21 1261 47
rect 1341 21 1371 47
rect 1425 21 1455 47
rect 1519 21 1549 47
rect 1613 21 1643 47
rect 1717 21 1747 47
rect 1801 21 1831 47
rect 1895 21 1925 47
rect 1989 21 2019 47
<< polycont >>
rect 81 215 115 249
rect 159 215 193 249
rect 237 215 271 249
rect 315 215 349 249
rect 570 215 604 249
rect 648 215 682 249
rect 726 215 760 249
rect 1035 215 1069 249
rect 1113 215 1147 249
rect 1219 215 1253 249
rect 1329 215 1363 249
rect 1519 215 1553 249
rect 1590 215 1624 249
rect 1675 215 1709 249
rect 1817 215 1851 249
rect 1895 215 1929 249
rect 1973 215 2007 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 31 483 81 527
rect 31 449 39 483
rect 73 449 81 483
rect 31 415 81 449
rect 31 381 39 415
rect 73 381 81 415
rect 31 347 81 381
rect 31 313 39 347
rect 73 313 81 347
rect 31 297 81 313
rect 125 477 175 493
rect 125 443 133 477
rect 167 443 175 477
rect 125 409 175 443
rect 125 375 133 409
rect 167 375 175 409
rect 125 341 175 375
rect 219 483 269 527
rect 219 449 227 483
rect 261 449 269 483
rect 219 415 269 449
rect 219 381 227 415
rect 261 381 269 415
rect 219 365 269 381
rect 313 477 363 493
rect 313 443 321 477
rect 355 443 363 477
rect 313 409 363 443
rect 407 477 561 527
rect 407 443 415 477
rect 449 443 519 477
rect 553 443 561 477
rect 407 425 561 443
rect 605 477 655 493
rect 605 443 613 477
rect 647 443 655 477
rect 313 375 321 409
rect 355 391 363 409
rect 605 409 655 443
rect 699 477 749 527
rect 699 443 707 477
rect 741 443 749 477
rect 699 425 749 443
rect 793 487 1227 493
rect 793 477 989 487
rect 793 443 801 477
rect 835 453 989 477
rect 1023 453 1177 487
rect 1211 453 1227 487
rect 1271 487 1321 527
rect 1271 453 1279 487
rect 1313 453 1321 487
rect 1355 487 1799 493
rect 1355 453 1381 487
rect 1415 453 1569 487
rect 1603 477 1799 487
rect 1603 453 1757 477
rect 355 375 465 391
rect 125 307 133 341
rect 167 323 175 341
rect 313 341 465 375
rect 605 375 613 409
rect 647 391 655 409
rect 793 409 835 443
rect 1271 435 1321 453
rect 1791 443 1799 477
rect 793 391 801 409
rect 647 375 801 391
rect 1757 409 1799 443
rect 1843 477 1893 527
rect 1843 443 1851 477
rect 1885 443 1893 477
rect 1843 425 1893 443
rect 1937 477 1987 493
rect 1937 443 1945 477
rect 1979 443 1987 477
rect 605 357 835 375
rect 869 367 895 401
rect 929 367 1083 401
rect 1117 367 1475 401
rect 1509 367 1663 401
rect 1697 367 1713 401
rect 869 357 1713 367
rect 1791 391 1799 409
rect 1937 409 1987 443
rect 1937 391 1945 409
rect 1791 375 1945 391
rect 1979 375 1987 409
rect 1757 357 1987 375
rect 313 323 321 341
rect 167 307 321 323
rect 355 323 465 341
rect 869 323 913 357
rect 1937 341 1987 357
rect 355 307 913 323
rect 125 289 913 307
rect 947 289 1279 323
rect 18 249 380 255
rect 18 215 81 249
rect 115 215 159 249
rect 193 215 237 249
rect 271 215 315 249
rect 349 215 380 249
rect 23 163 73 179
rect 424 173 465 289
rect 947 255 985 289
rect 512 249 985 255
rect 512 215 570 249
rect 604 215 648 249
rect 682 215 726 249
rect 760 215 985 249
rect 1019 249 1167 255
rect 1019 215 1035 249
rect 1069 215 1113 249
rect 1147 215 1167 249
rect 1203 249 1279 289
rect 1203 215 1219 249
rect 1253 215 1279 249
rect 1313 289 1864 323
rect 1937 307 1945 341
rect 1979 307 1987 341
rect 1937 289 1987 307
rect 2031 477 2081 527
rect 2031 443 2039 477
rect 2073 443 2081 477
rect 2031 409 2081 443
rect 2031 375 2039 409
rect 2073 375 2081 409
rect 2031 341 2081 375
rect 2031 307 2039 341
rect 2073 307 2081 341
rect 2031 289 2081 307
rect 1313 249 1389 289
rect 1801 255 1864 289
rect 1313 215 1329 249
rect 1363 215 1389 249
rect 1425 249 1747 255
rect 1425 215 1519 249
rect 1553 215 1590 249
rect 1624 215 1675 249
rect 1709 215 1747 249
rect 1801 249 2027 255
rect 1801 215 1817 249
rect 1851 215 1895 249
rect 1929 215 1973 249
rect 2007 215 2027 249
rect 1019 199 1167 215
rect 23 129 39 163
rect 107 163 465 173
rect 1203 164 2089 181
rect 107 129 133 163
rect 167 129 321 163
rect 355 129 465 163
rect 503 163 2089 164
rect 503 129 519 163
rect 553 129 707 163
rect 741 129 895 163
rect 929 129 1083 163
rect 1117 129 1287 163
rect 1321 147 1475 163
rect 1321 129 1337 147
rect 23 95 73 129
rect 1271 95 1337 129
rect 1449 129 1475 147
rect 1509 145 1663 163
rect 1509 129 1525 145
rect 23 61 39 95
rect 73 61 227 95
rect 261 61 415 95
rect 449 61 613 95
rect 647 61 801 95
rect 835 61 989 95
rect 1023 61 1177 95
rect 1211 61 1227 95
rect 23 51 1227 61
rect 1271 61 1287 95
rect 1321 61 1337 95
rect 1271 51 1337 61
rect 1381 95 1415 111
rect 1381 17 1415 61
rect 1449 95 1525 129
rect 1637 129 1663 145
rect 1697 147 1851 163
rect 1697 129 1713 147
rect 1449 61 1475 95
rect 1509 61 1525 95
rect 1449 51 1525 61
rect 1569 95 1603 111
rect 1569 17 1603 61
rect 1637 95 1713 129
rect 1825 129 1851 147
rect 1885 145 2039 163
rect 1885 129 1901 145
rect 1637 61 1663 95
rect 1697 61 1713 95
rect 1637 51 1713 61
rect 1757 95 1791 111
rect 1757 17 1791 61
rect 1825 95 1901 129
rect 2013 129 2039 145
rect 2073 129 2089 163
rect 1825 61 1851 95
rect 1885 61 1901 95
rect 1825 51 1901 61
rect 1945 95 1979 111
rect 1945 17 1979 61
rect 2013 95 2089 129
rect 2013 61 2039 95
rect 2073 61 2089 95
rect 2013 51 2089 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< labels >>
flabel locali s 1203 215 1279 289 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 1019 199 1167 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 1564 221 1598 255 0 FreeSans 400 180 0 0 A2
port 2 nsew signal input
flabel locali s 211 221 245 255 0 FreeSans 400 0 0 0 C1
port 5 nsew signal input
flabel locali s 1317 357 1351 391 0 FreeSans 400 180 0 0 Y
port 10 nsew signal output
flabel locali s 1870 221 1904 255 0 FreeSans 400 180 0 0 A1
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221ai_4
rlabel locali s 947 289 1279 323 1 B1
port 3 nsew signal input
rlabel locali s 947 255 985 289 1 B1
port 3 nsew signal input
rlabel locali s 512 215 985 255 1 B1
port 3 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 2116 544
string GDS_END 2041130
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 2027060
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
