magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 560 203
rect 29 -17 63 21
<< scnmos >>
rect 83 47 113 177
rect 272 47 302 177
rect 356 47 386 177
rect 452 47 482 177
<< scpmoshvt >>
rect 85 297 121 497
rect 250 297 286 497
rect 358 297 394 497
rect 454 297 490 497
<< ndiff >>
rect 27 164 83 177
rect 27 130 35 164
rect 69 130 83 164
rect 27 96 83 130
rect 27 62 35 96
rect 69 62 83 96
rect 27 47 83 62
rect 113 93 165 177
rect 113 59 123 93
rect 157 59 165 93
rect 113 47 165 59
rect 219 165 272 177
rect 219 131 227 165
rect 261 131 272 165
rect 219 97 272 131
rect 219 63 227 97
rect 261 63 272 97
rect 219 47 272 63
rect 302 161 356 177
rect 302 127 312 161
rect 346 127 356 161
rect 302 47 356 127
rect 386 93 452 177
rect 386 59 396 93
rect 430 59 452 93
rect 386 47 452 59
rect 482 165 534 177
rect 482 131 492 165
rect 526 131 534 165
rect 482 97 534 131
rect 482 63 492 97
rect 526 63 534 97
rect 482 47 534 63
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 485 250 497
rect 121 383 135 485
rect 237 383 250 485
rect 121 297 250 383
rect 286 485 358 497
rect 286 451 312 485
rect 346 451 358 485
rect 286 417 358 451
rect 286 383 312 417
rect 346 383 358 417
rect 286 349 358 383
rect 286 315 312 349
rect 346 315 358 349
rect 286 297 358 315
rect 394 297 454 497
rect 490 485 612 497
rect 490 383 502 485
rect 604 383 612 485
rect 490 297 612 383
<< ndiffc >>
rect 35 130 69 164
rect 35 62 69 96
rect 123 59 157 93
rect 227 131 261 165
rect 227 63 261 97
rect 312 127 346 161
rect 396 59 430 93
rect 492 131 526 165
rect 492 63 526 97
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 135 383 237 485
rect 312 451 346 485
rect 312 383 346 417
rect 312 315 346 349
rect 502 383 604 485
<< poly >>
rect 85 497 121 523
rect 250 497 286 523
rect 358 497 394 523
rect 454 497 490 523
rect 85 282 121 297
rect 250 282 286 297
rect 358 282 394 297
rect 454 282 490 297
rect 83 265 123 282
rect 248 265 288 282
rect 356 265 396 282
rect 452 269 492 282
rect 83 249 164 265
rect 83 215 120 249
rect 154 215 164 249
rect 83 199 164 215
rect 248 249 302 265
rect 248 215 258 249
rect 292 215 302 249
rect 248 199 302 215
rect 83 177 113 199
rect 272 177 302 199
rect 356 249 410 265
rect 356 215 366 249
rect 400 215 410 249
rect 356 199 410 215
rect 452 249 525 269
rect 452 215 481 249
rect 515 215 525 249
rect 452 199 525 215
rect 356 177 386 199
rect 452 177 482 199
rect 83 21 113 47
rect 272 21 302 47
rect 356 21 386 47
rect 452 21 482 47
<< polycont >>
rect 120 215 154 249
rect 258 215 292 249
rect 366 215 400 249
rect 481 215 515 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 477 73 493
rect 17 443 39 477
rect 17 409 73 443
rect 17 375 39 409
rect 17 341 73 375
rect 107 485 253 527
rect 107 383 135 485
rect 237 383 253 485
rect 107 372 253 383
rect 296 485 362 493
rect 296 451 312 485
rect 346 451 362 485
rect 476 485 620 527
rect 296 417 362 451
rect 296 383 312 417
rect 346 383 362 417
rect 17 307 39 341
rect 296 349 362 383
rect 296 338 312 349
rect 17 206 73 307
rect 120 315 312 338
rect 346 315 362 349
rect 120 295 362 315
rect 120 249 177 295
rect 154 215 177 249
rect 211 249 311 261
rect 397 255 431 478
rect 476 383 502 485
rect 604 383 620 485
rect 211 215 258 249
rect 292 215 311 249
rect 345 249 431 255
rect 345 215 366 249
rect 400 215 431 249
rect 465 249 535 323
rect 465 215 481 249
rect 515 215 535 249
rect 17 164 85 206
rect 17 130 35 164
rect 69 130 85 164
rect 120 181 177 215
rect 120 165 277 181
rect 120 143 227 165
rect 17 96 85 130
rect 205 131 227 143
rect 261 131 277 165
rect 17 62 35 96
rect 69 62 85 96
rect 17 51 85 62
rect 123 93 157 109
rect 123 17 157 59
rect 205 97 277 131
rect 311 165 542 181
rect 311 161 492 165
rect 311 127 312 161
rect 346 143 492 161
rect 346 127 353 143
rect 311 111 353 127
rect 476 131 492 143
rect 526 131 542 165
rect 205 63 227 97
rect 261 63 277 97
rect 205 51 277 63
rect 396 93 430 109
rect 396 17 430 59
rect 476 97 542 131
rect 476 63 492 97
rect 526 63 542 97
rect 476 51 542 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 29 357 63 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 465 289 499 323 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 211 215 311 261 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 364 221 398 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21a_1
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 1903126
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1897362
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
