magic
tech sky130A
magscale 1 2
timestamp 1729812420
<< metal3 >>
rect -892 11372 -120 11400
rect -892 10948 -204 11372
rect -140 10948 -120 11372
rect -892 10920 -120 10948
rect 120 11372 892 11400
rect 120 10948 808 11372
rect 872 10948 892 11372
rect 120 10920 892 10948
rect -892 10652 -120 10680
rect -892 10228 -204 10652
rect -140 10228 -120 10652
rect -892 10200 -120 10228
rect 120 10652 892 10680
rect 120 10228 808 10652
rect 872 10228 892 10652
rect 120 10200 892 10228
rect -892 9932 -120 9960
rect -892 9508 -204 9932
rect -140 9508 -120 9932
rect -892 9480 -120 9508
rect 120 9932 892 9960
rect 120 9508 808 9932
rect 872 9508 892 9932
rect 120 9480 892 9508
rect -892 9212 -120 9240
rect -892 8788 -204 9212
rect -140 8788 -120 9212
rect -892 8760 -120 8788
rect 120 9212 892 9240
rect 120 8788 808 9212
rect 872 8788 892 9212
rect 120 8760 892 8788
rect -892 8492 -120 8520
rect -892 8068 -204 8492
rect -140 8068 -120 8492
rect -892 8040 -120 8068
rect 120 8492 892 8520
rect 120 8068 808 8492
rect 872 8068 892 8492
rect 120 8040 892 8068
rect -892 7772 -120 7800
rect -892 7348 -204 7772
rect -140 7348 -120 7772
rect -892 7320 -120 7348
rect 120 7772 892 7800
rect 120 7348 808 7772
rect 872 7348 892 7772
rect 120 7320 892 7348
rect -892 7052 -120 7080
rect -892 6628 -204 7052
rect -140 6628 -120 7052
rect -892 6600 -120 6628
rect 120 7052 892 7080
rect 120 6628 808 7052
rect 872 6628 892 7052
rect 120 6600 892 6628
rect -892 6332 -120 6360
rect -892 5908 -204 6332
rect -140 5908 -120 6332
rect -892 5880 -120 5908
rect 120 6332 892 6360
rect 120 5908 808 6332
rect 872 5908 892 6332
rect 120 5880 892 5908
rect -892 5612 -120 5640
rect -892 5188 -204 5612
rect -140 5188 -120 5612
rect -892 5160 -120 5188
rect 120 5612 892 5640
rect 120 5188 808 5612
rect 872 5188 892 5612
rect 120 5160 892 5188
rect -892 4892 -120 4920
rect -892 4468 -204 4892
rect -140 4468 -120 4892
rect -892 4440 -120 4468
rect 120 4892 892 4920
rect 120 4468 808 4892
rect 872 4468 892 4892
rect 120 4440 892 4468
rect -892 4172 -120 4200
rect -892 3748 -204 4172
rect -140 3748 -120 4172
rect -892 3720 -120 3748
rect 120 4172 892 4200
rect 120 3748 808 4172
rect 872 3748 892 4172
rect 120 3720 892 3748
rect -892 3452 -120 3480
rect -892 3028 -204 3452
rect -140 3028 -120 3452
rect -892 3000 -120 3028
rect 120 3452 892 3480
rect 120 3028 808 3452
rect 872 3028 892 3452
rect 120 3000 892 3028
rect -892 2732 -120 2760
rect -892 2308 -204 2732
rect -140 2308 -120 2732
rect -892 2280 -120 2308
rect 120 2732 892 2760
rect 120 2308 808 2732
rect 872 2308 892 2732
rect 120 2280 892 2308
rect -892 2012 -120 2040
rect -892 1588 -204 2012
rect -140 1588 -120 2012
rect -892 1560 -120 1588
rect 120 2012 892 2040
rect 120 1588 808 2012
rect 872 1588 892 2012
rect 120 1560 892 1588
rect -892 1292 -120 1320
rect -892 868 -204 1292
rect -140 868 -120 1292
rect -892 840 -120 868
rect 120 1292 892 1320
rect 120 868 808 1292
rect 872 868 892 1292
rect 120 840 892 868
rect -892 572 -120 600
rect -892 148 -204 572
rect -140 148 -120 572
rect -892 120 -120 148
rect 120 572 892 600
rect 120 148 808 572
rect 872 148 892 572
rect 120 120 892 148
rect -892 -148 -120 -120
rect -892 -572 -204 -148
rect -140 -572 -120 -148
rect -892 -600 -120 -572
rect 120 -148 892 -120
rect 120 -572 808 -148
rect 872 -572 892 -148
rect 120 -600 892 -572
rect -892 -868 -120 -840
rect -892 -1292 -204 -868
rect -140 -1292 -120 -868
rect -892 -1320 -120 -1292
rect 120 -868 892 -840
rect 120 -1292 808 -868
rect 872 -1292 892 -868
rect 120 -1320 892 -1292
rect -892 -1588 -120 -1560
rect -892 -2012 -204 -1588
rect -140 -2012 -120 -1588
rect -892 -2040 -120 -2012
rect 120 -1588 892 -1560
rect 120 -2012 808 -1588
rect 872 -2012 892 -1588
rect 120 -2040 892 -2012
rect -892 -2308 -120 -2280
rect -892 -2732 -204 -2308
rect -140 -2732 -120 -2308
rect -892 -2760 -120 -2732
rect 120 -2308 892 -2280
rect 120 -2732 808 -2308
rect 872 -2732 892 -2308
rect 120 -2760 892 -2732
rect -892 -3028 -120 -3000
rect -892 -3452 -204 -3028
rect -140 -3452 -120 -3028
rect -892 -3480 -120 -3452
rect 120 -3028 892 -3000
rect 120 -3452 808 -3028
rect 872 -3452 892 -3028
rect 120 -3480 892 -3452
rect -892 -3748 -120 -3720
rect -892 -4172 -204 -3748
rect -140 -4172 -120 -3748
rect -892 -4200 -120 -4172
rect 120 -3748 892 -3720
rect 120 -4172 808 -3748
rect 872 -4172 892 -3748
rect 120 -4200 892 -4172
rect -892 -4468 -120 -4440
rect -892 -4892 -204 -4468
rect -140 -4892 -120 -4468
rect -892 -4920 -120 -4892
rect 120 -4468 892 -4440
rect 120 -4892 808 -4468
rect 872 -4892 892 -4468
rect 120 -4920 892 -4892
rect -892 -5188 -120 -5160
rect -892 -5612 -204 -5188
rect -140 -5612 -120 -5188
rect -892 -5640 -120 -5612
rect 120 -5188 892 -5160
rect 120 -5612 808 -5188
rect 872 -5612 892 -5188
rect 120 -5640 892 -5612
rect -892 -5908 -120 -5880
rect -892 -6332 -204 -5908
rect -140 -6332 -120 -5908
rect -892 -6360 -120 -6332
rect 120 -5908 892 -5880
rect 120 -6332 808 -5908
rect 872 -6332 892 -5908
rect 120 -6360 892 -6332
rect -892 -6628 -120 -6600
rect -892 -7052 -204 -6628
rect -140 -7052 -120 -6628
rect -892 -7080 -120 -7052
rect 120 -6628 892 -6600
rect 120 -7052 808 -6628
rect 872 -7052 892 -6628
rect 120 -7080 892 -7052
rect -892 -7348 -120 -7320
rect -892 -7772 -204 -7348
rect -140 -7772 -120 -7348
rect -892 -7800 -120 -7772
rect 120 -7348 892 -7320
rect 120 -7772 808 -7348
rect 872 -7772 892 -7348
rect 120 -7800 892 -7772
rect -892 -8068 -120 -8040
rect -892 -8492 -204 -8068
rect -140 -8492 -120 -8068
rect -892 -8520 -120 -8492
rect 120 -8068 892 -8040
rect 120 -8492 808 -8068
rect 872 -8492 892 -8068
rect 120 -8520 892 -8492
rect -892 -8788 -120 -8760
rect -892 -9212 -204 -8788
rect -140 -9212 -120 -8788
rect -892 -9240 -120 -9212
rect 120 -8788 892 -8760
rect 120 -9212 808 -8788
rect 872 -9212 892 -8788
rect 120 -9240 892 -9212
rect -892 -9508 -120 -9480
rect -892 -9932 -204 -9508
rect -140 -9932 -120 -9508
rect -892 -9960 -120 -9932
rect 120 -9508 892 -9480
rect 120 -9932 808 -9508
rect 872 -9932 892 -9508
rect 120 -9960 892 -9932
rect -892 -10228 -120 -10200
rect -892 -10652 -204 -10228
rect -140 -10652 -120 -10228
rect -892 -10680 -120 -10652
rect 120 -10228 892 -10200
rect 120 -10652 808 -10228
rect 872 -10652 892 -10228
rect 120 -10680 892 -10652
rect -892 -10948 -120 -10920
rect -892 -11372 -204 -10948
rect -140 -11372 -120 -10948
rect -892 -11400 -120 -11372
rect 120 -10948 892 -10920
rect 120 -11372 808 -10948
rect 872 -11372 892 -10948
rect 120 -11400 892 -11372
<< via3 >>
rect -204 10948 -140 11372
rect 808 10948 872 11372
rect -204 10228 -140 10652
rect 808 10228 872 10652
rect -204 9508 -140 9932
rect 808 9508 872 9932
rect -204 8788 -140 9212
rect 808 8788 872 9212
rect -204 8068 -140 8492
rect 808 8068 872 8492
rect -204 7348 -140 7772
rect 808 7348 872 7772
rect -204 6628 -140 7052
rect 808 6628 872 7052
rect -204 5908 -140 6332
rect 808 5908 872 6332
rect -204 5188 -140 5612
rect 808 5188 872 5612
rect -204 4468 -140 4892
rect 808 4468 872 4892
rect -204 3748 -140 4172
rect 808 3748 872 4172
rect -204 3028 -140 3452
rect 808 3028 872 3452
rect -204 2308 -140 2732
rect 808 2308 872 2732
rect -204 1588 -140 2012
rect 808 1588 872 2012
rect -204 868 -140 1292
rect 808 868 872 1292
rect -204 148 -140 572
rect 808 148 872 572
rect -204 -572 -140 -148
rect 808 -572 872 -148
rect -204 -1292 -140 -868
rect 808 -1292 872 -868
rect -204 -2012 -140 -1588
rect 808 -2012 872 -1588
rect -204 -2732 -140 -2308
rect 808 -2732 872 -2308
rect -204 -3452 -140 -3028
rect 808 -3452 872 -3028
rect -204 -4172 -140 -3748
rect 808 -4172 872 -3748
rect -204 -4892 -140 -4468
rect 808 -4892 872 -4468
rect -204 -5612 -140 -5188
rect 808 -5612 872 -5188
rect -204 -6332 -140 -5908
rect 808 -6332 872 -5908
rect -204 -7052 -140 -6628
rect 808 -7052 872 -6628
rect -204 -7772 -140 -7348
rect 808 -7772 872 -7348
rect -204 -8492 -140 -8068
rect 808 -8492 872 -8068
rect -204 -9212 -140 -8788
rect 808 -9212 872 -8788
rect -204 -9932 -140 -9508
rect 808 -9932 872 -9508
rect -204 -10652 -140 -10228
rect 808 -10652 872 -10228
rect -204 -11372 -140 -10948
rect 808 -11372 872 -10948
<< mimcap >>
rect -852 11320 -452 11360
rect -852 11000 -812 11320
rect -492 11000 -452 11320
rect -852 10960 -452 11000
rect 160 11320 560 11360
rect 160 11000 200 11320
rect 520 11000 560 11320
rect 160 10960 560 11000
rect -852 10600 -452 10640
rect -852 10280 -812 10600
rect -492 10280 -452 10600
rect -852 10240 -452 10280
rect 160 10600 560 10640
rect 160 10280 200 10600
rect 520 10280 560 10600
rect 160 10240 560 10280
rect -852 9880 -452 9920
rect -852 9560 -812 9880
rect -492 9560 -452 9880
rect -852 9520 -452 9560
rect 160 9880 560 9920
rect 160 9560 200 9880
rect 520 9560 560 9880
rect 160 9520 560 9560
rect -852 9160 -452 9200
rect -852 8840 -812 9160
rect -492 8840 -452 9160
rect -852 8800 -452 8840
rect 160 9160 560 9200
rect 160 8840 200 9160
rect 520 8840 560 9160
rect 160 8800 560 8840
rect -852 8440 -452 8480
rect -852 8120 -812 8440
rect -492 8120 -452 8440
rect -852 8080 -452 8120
rect 160 8440 560 8480
rect 160 8120 200 8440
rect 520 8120 560 8440
rect 160 8080 560 8120
rect -852 7720 -452 7760
rect -852 7400 -812 7720
rect -492 7400 -452 7720
rect -852 7360 -452 7400
rect 160 7720 560 7760
rect 160 7400 200 7720
rect 520 7400 560 7720
rect 160 7360 560 7400
rect -852 7000 -452 7040
rect -852 6680 -812 7000
rect -492 6680 -452 7000
rect -852 6640 -452 6680
rect 160 7000 560 7040
rect 160 6680 200 7000
rect 520 6680 560 7000
rect 160 6640 560 6680
rect -852 6280 -452 6320
rect -852 5960 -812 6280
rect -492 5960 -452 6280
rect -852 5920 -452 5960
rect 160 6280 560 6320
rect 160 5960 200 6280
rect 520 5960 560 6280
rect 160 5920 560 5960
rect -852 5560 -452 5600
rect -852 5240 -812 5560
rect -492 5240 -452 5560
rect -852 5200 -452 5240
rect 160 5560 560 5600
rect 160 5240 200 5560
rect 520 5240 560 5560
rect 160 5200 560 5240
rect -852 4840 -452 4880
rect -852 4520 -812 4840
rect -492 4520 -452 4840
rect -852 4480 -452 4520
rect 160 4840 560 4880
rect 160 4520 200 4840
rect 520 4520 560 4840
rect 160 4480 560 4520
rect -852 4120 -452 4160
rect -852 3800 -812 4120
rect -492 3800 -452 4120
rect -852 3760 -452 3800
rect 160 4120 560 4160
rect 160 3800 200 4120
rect 520 3800 560 4120
rect 160 3760 560 3800
rect -852 3400 -452 3440
rect -852 3080 -812 3400
rect -492 3080 -452 3400
rect -852 3040 -452 3080
rect 160 3400 560 3440
rect 160 3080 200 3400
rect 520 3080 560 3400
rect 160 3040 560 3080
rect -852 2680 -452 2720
rect -852 2360 -812 2680
rect -492 2360 -452 2680
rect -852 2320 -452 2360
rect 160 2680 560 2720
rect 160 2360 200 2680
rect 520 2360 560 2680
rect 160 2320 560 2360
rect -852 1960 -452 2000
rect -852 1640 -812 1960
rect -492 1640 -452 1960
rect -852 1600 -452 1640
rect 160 1960 560 2000
rect 160 1640 200 1960
rect 520 1640 560 1960
rect 160 1600 560 1640
rect -852 1240 -452 1280
rect -852 920 -812 1240
rect -492 920 -452 1240
rect -852 880 -452 920
rect 160 1240 560 1280
rect 160 920 200 1240
rect 520 920 560 1240
rect 160 880 560 920
rect -852 520 -452 560
rect -852 200 -812 520
rect -492 200 -452 520
rect -852 160 -452 200
rect 160 520 560 560
rect 160 200 200 520
rect 520 200 560 520
rect 160 160 560 200
rect -852 -200 -452 -160
rect -852 -520 -812 -200
rect -492 -520 -452 -200
rect -852 -560 -452 -520
rect 160 -200 560 -160
rect 160 -520 200 -200
rect 520 -520 560 -200
rect 160 -560 560 -520
rect -852 -920 -452 -880
rect -852 -1240 -812 -920
rect -492 -1240 -452 -920
rect -852 -1280 -452 -1240
rect 160 -920 560 -880
rect 160 -1240 200 -920
rect 520 -1240 560 -920
rect 160 -1280 560 -1240
rect -852 -1640 -452 -1600
rect -852 -1960 -812 -1640
rect -492 -1960 -452 -1640
rect -852 -2000 -452 -1960
rect 160 -1640 560 -1600
rect 160 -1960 200 -1640
rect 520 -1960 560 -1640
rect 160 -2000 560 -1960
rect -852 -2360 -452 -2320
rect -852 -2680 -812 -2360
rect -492 -2680 -452 -2360
rect -852 -2720 -452 -2680
rect 160 -2360 560 -2320
rect 160 -2680 200 -2360
rect 520 -2680 560 -2360
rect 160 -2720 560 -2680
rect -852 -3080 -452 -3040
rect -852 -3400 -812 -3080
rect -492 -3400 -452 -3080
rect -852 -3440 -452 -3400
rect 160 -3080 560 -3040
rect 160 -3400 200 -3080
rect 520 -3400 560 -3080
rect 160 -3440 560 -3400
rect -852 -3800 -452 -3760
rect -852 -4120 -812 -3800
rect -492 -4120 -452 -3800
rect -852 -4160 -452 -4120
rect 160 -3800 560 -3760
rect 160 -4120 200 -3800
rect 520 -4120 560 -3800
rect 160 -4160 560 -4120
rect -852 -4520 -452 -4480
rect -852 -4840 -812 -4520
rect -492 -4840 -452 -4520
rect -852 -4880 -452 -4840
rect 160 -4520 560 -4480
rect 160 -4840 200 -4520
rect 520 -4840 560 -4520
rect 160 -4880 560 -4840
rect -852 -5240 -452 -5200
rect -852 -5560 -812 -5240
rect -492 -5560 -452 -5240
rect -852 -5600 -452 -5560
rect 160 -5240 560 -5200
rect 160 -5560 200 -5240
rect 520 -5560 560 -5240
rect 160 -5600 560 -5560
rect -852 -5960 -452 -5920
rect -852 -6280 -812 -5960
rect -492 -6280 -452 -5960
rect -852 -6320 -452 -6280
rect 160 -5960 560 -5920
rect 160 -6280 200 -5960
rect 520 -6280 560 -5960
rect 160 -6320 560 -6280
rect -852 -6680 -452 -6640
rect -852 -7000 -812 -6680
rect -492 -7000 -452 -6680
rect -852 -7040 -452 -7000
rect 160 -6680 560 -6640
rect 160 -7000 200 -6680
rect 520 -7000 560 -6680
rect 160 -7040 560 -7000
rect -852 -7400 -452 -7360
rect -852 -7720 -812 -7400
rect -492 -7720 -452 -7400
rect -852 -7760 -452 -7720
rect 160 -7400 560 -7360
rect 160 -7720 200 -7400
rect 520 -7720 560 -7400
rect 160 -7760 560 -7720
rect -852 -8120 -452 -8080
rect -852 -8440 -812 -8120
rect -492 -8440 -452 -8120
rect -852 -8480 -452 -8440
rect 160 -8120 560 -8080
rect 160 -8440 200 -8120
rect 520 -8440 560 -8120
rect 160 -8480 560 -8440
rect -852 -8840 -452 -8800
rect -852 -9160 -812 -8840
rect -492 -9160 -452 -8840
rect -852 -9200 -452 -9160
rect 160 -8840 560 -8800
rect 160 -9160 200 -8840
rect 520 -9160 560 -8840
rect 160 -9200 560 -9160
rect -852 -9560 -452 -9520
rect -852 -9880 -812 -9560
rect -492 -9880 -452 -9560
rect -852 -9920 -452 -9880
rect 160 -9560 560 -9520
rect 160 -9880 200 -9560
rect 520 -9880 560 -9560
rect 160 -9920 560 -9880
rect -852 -10280 -452 -10240
rect -852 -10600 -812 -10280
rect -492 -10600 -452 -10280
rect -852 -10640 -452 -10600
rect 160 -10280 560 -10240
rect 160 -10600 200 -10280
rect 520 -10600 560 -10280
rect 160 -10640 560 -10600
rect -852 -11000 -452 -10960
rect -852 -11320 -812 -11000
rect -492 -11320 -452 -11000
rect -852 -11360 -452 -11320
rect 160 -11000 560 -10960
rect 160 -11320 200 -11000
rect 520 -11320 560 -11000
rect 160 -11360 560 -11320
<< mimcapcontact >>
rect -812 11000 -492 11320
rect 200 11000 520 11320
rect -812 10280 -492 10600
rect 200 10280 520 10600
rect -812 9560 -492 9880
rect 200 9560 520 9880
rect -812 8840 -492 9160
rect 200 8840 520 9160
rect -812 8120 -492 8440
rect 200 8120 520 8440
rect -812 7400 -492 7720
rect 200 7400 520 7720
rect -812 6680 -492 7000
rect 200 6680 520 7000
rect -812 5960 -492 6280
rect 200 5960 520 6280
rect -812 5240 -492 5560
rect 200 5240 520 5560
rect -812 4520 -492 4840
rect 200 4520 520 4840
rect -812 3800 -492 4120
rect 200 3800 520 4120
rect -812 3080 -492 3400
rect 200 3080 520 3400
rect -812 2360 -492 2680
rect 200 2360 520 2680
rect -812 1640 -492 1960
rect 200 1640 520 1960
rect -812 920 -492 1240
rect 200 920 520 1240
rect -812 200 -492 520
rect 200 200 520 520
rect -812 -520 -492 -200
rect 200 -520 520 -200
rect -812 -1240 -492 -920
rect 200 -1240 520 -920
rect -812 -1960 -492 -1640
rect 200 -1960 520 -1640
rect -812 -2680 -492 -2360
rect 200 -2680 520 -2360
rect -812 -3400 -492 -3080
rect 200 -3400 520 -3080
rect -812 -4120 -492 -3800
rect 200 -4120 520 -3800
rect -812 -4840 -492 -4520
rect 200 -4840 520 -4520
rect -812 -5560 -492 -5240
rect 200 -5560 520 -5240
rect -812 -6280 -492 -5960
rect 200 -6280 520 -5960
rect -812 -7000 -492 -6680
rect 200 -7000 520 -6680
rect -812 -7720 -492 -7400
rect 200 -7720 520 -7400
rect -812 -8440 -492 -8120
rect 200 -8440 520 -8120
rect -812 -9160 -492 -8840
rect 200 -9160 520 -8840
rect -812 -9880 -492 -9560
rect 200 -9880 520 -9560
rect -812 -10600 -492 -10280
rect 200 -10600 520 -10280
rect -812 -11320 -492 -11000
rect 200 -11320 520 -11000
<< metal4 >>
rect -704 11321 -600 11520
rect -220 11372 -124 11388
rect -813 11320 -491 11321
rect -813 11000 -812 11320
rect -492 11000 -491 11320
rect -813 10999 -491 11000
rect -704 10601 -600 10999
rect -220 10948 -204 11372
rect -140 10948 -124 11372
rect 308 11321 412 11520
rect 792 11372 888 11388
rect 199 11320 521 11321
rect 199 11000 200 11320
rect 520 11000 521 11320
rect 199 10999 521 11000
rect -220 10932 -124 10948
rect -220 10652 -124 10668
rect -813 10600 -491 10601
rect -813 10280 -812 10600
rect -492 10280 -491 10600
rect -813 10279 -491 10280
rect -704 9881 -600 10279
rect -220 10228 -204 10652
rect -140 10228 -124 10652
rect 308 10601 412 10999
rect 792 10948 808 11372
rect 872 10948 888 11372
rect 792 10932 888 10948
rect 792 10652 888 10668
rect 199 10600 521 10601
rect 199 10280 200 10600
rect 520 10280 521 10600
rect 199 10279 521 10280
rect -220 10212 -124 10228
rect -220 9932 -124 9948
rect -813 9880 -491 9881
rect -813 9560 -812 9880
rect -492 9560 -491 9880
rect -813 9559 -491 9560
rect -704 9161 -600 9559
rect -220 9508 -204 9932
rect -140 9508 -124 9932
rect 308 9881 412 10279
rect 792 10228 808 10652
rect 872 10228 888 10652
rect 792 10212 888 10228
rect 792 9932 888 9948
rect 199 9880 521 9881
rect 199 9560 200 9880
rect 520 9560 521 9880
rect 199 9559 521 9560
rect -220 9492 -124 9508
rect -220 9212 -124 9228
rect -813 9160 -491 9161
rect -813 8840 -812 9160
rect -492 8840 -491 9160
rect -813 8839 -491 8840
rect -704 8441 -600 8839
rect -220 8788 -204 9212
rect -140 8788 -124 9212
rect 308 9161 412 9559
rect 792 9508 808 9932
rect 872 9508 888 9932
rect 792 9492 888 9508
rect 792 9212 888 9228
rect 199 9160 521 9161
rect 199 8840 200 9160
rect 520 8840 521 9160
rect 199 8839 521 8840
rect -220 8772 -124 8788
rect -220 8492 -124 8508
rect -813 8440 -491 8441
rect -813 8120 -812 8440
rect -492 8120 -491 8440
rect -813 8119 -491 8120
rect -704 7721 -600 8119
rect -220 8068 -204 8492
rect -140 8068 -124 8492
rect 308 8441 412 8839
rect 792 8788 808 9212
rect 872 8788 888 9212
rect 792 8772 888 8788
rect 792 8492 888 8508
rect 199 8440 521 8441
rect 199 8120 200 8440
rect 520 8120 521 8440
rect 199 8119 521 8120
rect -220 8052 -124 8068
rect -220 7772 -124 7788
rect -813 7720 -491 7721
rect -813 7400 -812 7720
rect -492 7400 -491 7720
rect -813 7399 -491 7400
rect -704 7001 -600 7399
rect -220 7348 -204 7772
rect -140 7348 -124 7772
rect 308 7721 412 8119
rect 792 8068 808 8492
rect 872 8068 888 8492
rect 792 8052 888 8068
rect 792 7772 888 7788
rect 199 7720 521 7721
rect 199 7400 200 7720
rect 520 7400 521 7720
rect 199 7399 521 7400
rect -220 7332 -124 7348
rect -220 7052 -124 7068
rect -813 7000 -491 7001
rect -813 6680 -812 7000
rect -492 6680 -491 7000
rect -813 6679 -491 6680
rect -704 6281 -600 6679
rect -220 6628 -204 7052
rect -140 6628 -124 7052
rect 308 7001 412 7399
rect 792 7348 808 7772
rect 872 7348 888 7772
rect 792 7332 888 7348
rect 792 7052 888 7068
rect 199 7000 521 7001
rect 199 6680 200 7000
rect 520 6680 521 7000
rect 199 6679 521 6680
rect -220 6612 -124 6628
rect -220 6332 -124 6348
rect -813 6280 -491 6281
rect -813 5960 -812 6280
rect -492 5960 -491 6280
rect -813 5959 -491 5960
rect -704 5561 -600 5959
rect -220 5908 -204 6332
rect -140 5908 -124 6332
rect 308 6281 412 6679
rect 792 6628 808 7052
rect 872 6628 888 7052
rect 792 6612 888 6628
rect 792 6332 888 6348
rect 199 6280 521 6281
rect 199 5960 200 6280
rect 520 5960 521 6280
rect 199 5959 521 5960
rect -220 5892 -124 5908
rect -220 5612 -124 5628
rect -813 5560 -491 5561
rect -813 5240 -812 5560
rect -492 5240 -491 5560
rect -813 5239 -491 5240
rect -704 4841 -600 5239
rect -220 5188 -204 5612
rect -140 5188 -124 5612
rect 308 5561 412 5959
rect 792 5908 808 6332
rect 872 5908 888 6332
rect 792 5892 888 5908
rect 792 5612 888 5628
rect 199 5560 521 5561
rect 199 5240 200 5560
rect 520 5240 521 5560
rect 199 5239 521 5240
rect -220 5172 -124 5188
rect -220 4892 -124 4908
rect -813 4840 -491 4841
rect -813 4520 -812 4840
rect -492 4520 -491 4840
rect -813 4519 -491 4520
rect -704 4121 -600 4519
rect -220 4468 -204 4892
rect -140 4468 -124 4892
rect 308 4841 412 5239
rect 792 5188 808 5612
rect 872 5188 888 5612
rect 792 5172 888 5188
rect 792 4892 888 4908
rect 199 4840 521 4841
rect 199 4520 200 4840
rect 520 4520 521 4840
rect 199 4519 521 4520
rect -220 4452 -124 4468
rect -220 4172 -124 4188
rect -813 4120 -491 4121
rect -813 3800 -812 4120
rect -492 3800 -491 4120
rect -813 3799 -491 3800
rect -704 3401 -600 3799
rect -220 3748 -204 4172
rect -140 3748 -124 4172
rect 308 4121 412 4519
rect 792 4468 808 4892
rect 872 4468 888 4892
rect 792 4452 888 4468
rect 792 4172 888 4188
rect 199 4120 521 4121
rect 199 3800 200 4120
rect 520 3800 521 4120
rect 199 3799 521 3800
rect -220 3732 -124 3748
rect -220 3452 -124 3468
rect -813 3400 -491 3401
rect -813 3080 -812 3400
rect -492 3080 -491 3400
rect -813 3079 -491 3080
rect -704 2681 -600 3079
rect -220 3028 -204 3452
rect -140 3028 -124 3452
rect 308 3401 412 3799
rect 792 3748 808 4172
rect 872 3748 888 4172
rect 792 3732 888 3748
rect 792 3452 888 3468
rect 199 3400 521 3401
rect 199 3080 200 3400
rect 520 3080 521 3400
rect 199 3079 521 3080
rect -220 3012 -124 3028
rect -220 2732 -124 2748
rect -813 2680 -491 2681
rect -813 2360 -812 2680
rect -492 2360 -491 2680
rect -813 2359 -491 2360
rect -704 1961 -600 2359
rect -220 2308 -204 2732
rect -140 2308 -124 2732
rect 308 2681 412 3079
rect 792 3028 808 3452
rect 872 3028 888 3452
rect 792 3012 888 3028
rect 792 2732 888 2748
rect 199 2680 521 2681
rect 199 2360 200 2680
rect 520 2360 521 2680
rect 199 2359 521 2360
rect -220 2292 -124 2308
rect -220 2012 -124 2028
rect -813 1960 -491 1961
rect -813 1640 -812 1960
rect -492 1640 -491 1960
rect -813 1639 -491 1640
rect -704 1241 -600 1639
rect -220 1588 -204 2012
rect -140 1588 -124 2012
rect 308 1961 412 2359
rect 792 2308 808 2732
rect 872 2308 888 2732
rect 792 2292 888 2308
rect 792 2012 888 2028
rect 199 1960 521 1961
rect 199 1640 200 1960
rect 520 1640 521 1960
rect 199 1639 521 1640
rect -220 1572 -124 1588
rect -220 1292 -124 1308
rect -813 1240 -491 1241
rect -813 920 -812 1240
rect -492 920 -491 1240
rect -813 919 -491 920
rect -704 521 -600 919
rect -220 868 -204 1292
rect -140 868 -124 1292
rect 308 1241 412 1639
rect 792 1588 808 2012
rect 872 1588 888 2012
rect 792 1572 888 1588
rect 792 1292 888 1308
rect 199 1240 521 1241
rect 199 920 200 1240
rect 520 920 521 1240
rect 199 919 521 920
rect -220 852 -124 868
rect -220 572 -124 588
rect -813 520 -491 521
rect -813 200 -812 520
rect -492 200 -491 520
rect -813 199 -491 200
rect -704 -199 -600 199
rect -220 148 -204 572
rect -140 148 -124 572
rect 308 521 412 919
rect 792 868 808 1292
rect 872 868 888 1292
rect 792 852 888 868
rect 792 572 888 588
rect 199 520 521 521
rect 199 200 200 520
rect 520 200 521 520
rect 199 199 521 200
rect -220 132 -124 148
rect -220 -148 -124 -132
rect -813 -200 -491 -199
rect -813 -520 -812 -200
rect -492 -520 -491 -200
rect -813 -521 -491 -520
rect -704 -919 -600 -521
rect -220 -572 -204 -148
rect -140 -572 -124 -148
rect 308 -199 412 199
rect 792 148 808 572
rect 872 148 888 572
rect 792 132 888 148
rect 792 -148 888 -132
rect 199 -200 521 -199
rect 199 -520 200 -200
rect 520 -520 521 -200
rect 199 -521 521 -520
rect -220 -588 -124 -572
rect -220 -868 -124 -852
rect -813 -920 -491 -919
rect -813 -1240 -812 -920
rect -492 -1240 -491 -920
rect -813 -1241 -491 -1240
rect -704 -1639 -600 -1241
rect -220 -1292 -204 -868
rect -140 -1292 -124 -868
rect 308 -919 412 -521
rect 792 -572 808 -148
rect 872 -572 888 -148
rect 792 -588 888 -572
rect 792 -868 888 -852
rect 199 -920 521 -919
rect 199 -1240 200 -920
rect 520 -1240 521 -920
rect 199 -1241 521 -1240
rect -220 -1308 -124 -1292
rect -220 -1588 -124 -1572
rect -813 -1640 -491 -1639
rect -813 -1960 -812 -1640
rect -492 -1960 -491 -1640
rect -813 -1961 -491 -1960
rect -704 -2359 -600 -1961
rect -220 -2012 -204 -1588
rect -140 -2012 -124 -1588
rect 308 -1639 412 -1241
rect 792 -1292 808 -868
rect 872 -1292 888 -868
rect 792 -1308 888 -1292
rect 792 -1588 888 -1572
rect 199 -1640 521 -1639
rect 199 -1960 200 -1640
rect 520 -1960 521 -1640
rect 199 -1961 521 -1960
rect -220 -2028 -124 -2012
rect -220 -2308 -124 -2292
rect -813 -2360 -491 -2359
rect -813 -2680 -812 -2360
rect -492 -2680 -491 -2360
rect -813 -2681 -491 -2680
rect -704 -3079 -600 -2681
rect -220 -2732 -204 -2308
rect -140 -2732 -124 -2308
rect 308 -2359 412 -1961
rect 792 -2012 808 -1588
rect 872 -2012 888 -1588
rect 792 -2028 888 -2012
rect 792 -2308 888 -2292
rect 199 -2360 521 -2359
rect 199 -2680 200 -2360
rect 520 -2680 521 -2360
rect 199 -2681 521 -2680
rect -220 -2748 -124 -2732
rect -220 -3028 -124 -3012
rect -813 -3080 -491 -3079
rect -813 -3400 -812 -3080
rect -492 -3400 -491 -3080
rect -813 -3401 -491 -3400
rect -704 -3799 -600 -3401
rect -220 -3452 -204 -3028
rect -140 -3452 -124 -3028
rect 308 -3079 412 -2681
rect 792 -2732 808 -2308
rect 872 -2732 888 -2308
rect 792 -2748 888 -2732
rect 792 -3028 888 -3012
rect 199 -3080 521 -3079
rect 199 -3400 200 -3080
rect 520 -3400 521 -3080
rect 199 -3401 521 -3400
rect -220 -3468 -124 -3452
rect -220 -3748 -124 -3732
rect -813 -3800 -491 -3799
rect -813 -4120 -812 -3800
rect -492 -4120 -491 -3800
rect -813 -4121 -491 -4120
rect -704 -4519 -600 -4121
rect -220 -4172 -204 -3748
rect -140 -4172 -124 -3748
rect 308 -3799 412 -3401
rect 792 -3452 808 -3028
rect 872 -3452 888 -3028
rect 792 -3468 888 -3452
rect 792 -3748 888 -3732
rect 199 -3800 521 -3799
rect 199 -4120 200 -3800
rect 520 -4120 521 -3800
rect 199 -4121 521 -4120
rect -220 -4188 -124 -4172
rect -220 -4468 -124 -4452
rect -813 -4520 -491 -4519
rect -813 -4840 -812 -4520
rect -492 -4840 -491 -4520
rect -813 -4841 -491 -4840
rect -704 -5239 -600 -4841
rect -220 -4892 -204 -4468
rect -140 -4892 -124 -4468
rect 308 -4519 412 -4121
rect 792 -4172 808 -3748
rect 872 -4172 888 -3748
rect 792 -4188 888 -4172
rect 792 -4468 888 -4452
rect 199 -4520 521 -4519
rect 199 -4840 200 -4520
rect 520 -4840 521 -4520
rect 199 -4841 521 -4840
rect -220 -4908 -124 -4892
rect -220 -5188 -124 -5172
rect -813 -5240 -491 -5239
rect -813 -5560 -812 -5240
rect -492 -5560 -491 -5240
rect -813 -5561 -491 -5560
rect -704 -5959 -600 -5561
rect -220 -5612 -204 -5188
rect -140 -5612 -124 -5188
rect 308 -5239 412 -4841
rect 792 -4892 808 -4468
rect 872 -4892 888 -4468
rect 792 -4908 888 -4892
rect 792 -5188 888 -5172
rect 199 -5240 521 -5239
rect 199 -5560 200 -5240
rect 520 -5560 521 -5240
rect 199 -5561 521 -5560
rect -220 -5628 -124 -5612
rect -220 -5908 -124 -5892
rect -813 -5960 -491 -5959
rect -813 -6280 -812 -5960
rect -492 -6280 -491 -5960
rect -813 -6281 -491 -6280
rect -704 -6679 -600 -6281
rect -220 -6332 -204 -5908
rect -140 -6332 -124 -5908
rect 308 -5959 412 -5561
rect 792 -5612 808 -5188
rect 872 -5612 888 -5188
rect 792 -5628 888 -5612
rect 792 -5908 888 -5892
rect 199 -5960 521 -5959
rect 199 -6280 200 -5960
rect 520 -6280 521 -5960
rect 199 -6281 521 -6280
rect -220 -6348 -124 -6332
rect -220 -6628 -124 -6612
rect -813 -6680 -491 -6679
rect -813 -7000 -812 -6680
rect -492 -7000 -491 -6680
rect -813 -7001 -491 -7000
rect -704 -7399 -600 -7001
rect -220 -7052 -204 -6628
rect -140 -7052 -124 -6628
rect 308 -6679 412 -6281
rect 792 -6332 808 -5908
rect 872 -6332 888 -5908
rect 792 -6348 888 -6332
rect 792 -6628 888 -6612
rect 199 -6680 521 -6679
rect 199 -7000 200 -6680
rect 520 -7000 521 -6680
rect 199 -7001 521 -7000
rect -220 -7068 -124 -7052
rect -220 -7348 -124 -7332
rect -813 -7400 -491 -7399
rect -813 -7720 -812 -7400
rect -492 -7720 -491 -7400
rect -813 -7721 -491 -7720
rect -704 -8119 -600 -7721
rect -220 -7772 -204 -7348
rect -140 -7772 -124 -7348
rect 308 -7399 412 -7001
rect 792 -7052 808 -6628
rect 872 -7052 888 -6628
rect 792 -7068 888 -7052
rect 792 -7348 888 -7332
rect 199 -7400 521 -7399
rect 199 -7720 200 -7400
rect 520 -7720 521 -7400
rect 199 -7721 521 -7720
rect -220 -7788 -124 -7772
rect -220 -8068 -124 -8052
rect -813 -8120 -491 -8119
rect -813 -8440 -812 -8120
rect -492 -8440 -491 -8120
rect -813 -8441 -491 -8440
rect -704 -8839 -600 -8441
rect -220 -8492 -204 -8068
rect -140 -8492 -124 -8068
rect 308 -8119 412 -7721
rect 792 -7772 808 -7348
rect 872 -7772 888 -7348
rect 792 -7788 888 -7772
rect 792 -8068 888 -8052
rect 199 -8120 521 -8119
rect 199 -8440 200 -8120
rect 520 -8440 521 -8120
rect 199 -8441 521 -8440
rect -220 -8508 -124 -8492
rect -220 -8788 -124 -8772
rect -813 -8840 -491 -8839
rect -813 -9160 -812 -8840
rect -492 -9160 -491 -8840
rect -813 -9161 -491 -9160
rect -704 -9559 -600 -9161
rect -220 -9212 -204 -8788
rect -140 -9212 -124 -8788
rect 308 -8839 412 -8441
rect 792 -8492 808 -8068
rect 872 -8492 888 -8068
rect 792 -8508 888 -8492
rect 792 -8788 888 -8772
rect 199 -8840 521 -8839
rect 199 -9160 200 -8840
rect 520 -9160 521 -8840
rect 199 -9161 521 -9160
rect -220 -9228 -124 -9212
rect -220 -9508 -124 -9492
rect -813 -9560 -491 -9559
rect -813 -9880 -812 -9560
rect -492 -9880 -491 -9560
rect -813 -9881 -491 -9880
rect -704 -10279 -600 -9881
rect -220 -9932 -204 -9508
rect -140 -9932 -124 -9508
rect 308 -9559 412 -9161
rect 792 -9212 808 -8788
rect 872 -9212 888 -8788
rect 792 -9228 888 -9212
rect 792 -9508 888 -9492
rect 199 -9560 521 -9559
rect 199 -9880 200 -9560
rect 520 -9880 521 -9560
rect 199 -9881 521 -9880
rect -220 -9948 -124 -9932
rect -220 -10228 -124 -10212
rect -813 -10280 -491 -10279
rect -813 -10600 -812 -10280
rect -492 -10600 -491 -10280
rect -813 -10601 -491 -10600
rect -704 -10999 -600 -10601
rect -220 -10652 -204 -10228
rect -140 -10652 -124 -10228
rect 308 -10279 412 -9881
rect 792 -9932 808 -9508
rect 872 -9932 888 -9508
rect 792 -9948 888 -9932
rect 792 -10228 888 -10212
rect 199 -10280 521 -10279
rect 199 -10600 200 -10280
rect 520 -10600 521 -10280
rect 199 -10601 521 -10600
rect -220 -10668 -124 -10652
rect -220 -10948 -124 -10932
rect -813 -11000 -491 -10999
rect -813 -11320 -812 -11000
rect -492 -11320 -491 -11000
rect -813 -11321 -491 -11320
rect -704 -11520 -600 -11321
rect -220 -11372 -204 -10948
rect -140 -11372 -124 -10948
rect 308 -10999 412 -10601
rect 792 -10652 808 -10228
rect 872 -10652 888 -10228
rect 792 -10668 888 -10652
rect 792 -10948 888 -10932
rect 199 -11000 521 -10999
rect 199 -11320 200 -11000
rect 520 -11320 521 -11000
rect 199 -11321 521 -11320
rect -220 -11388 -124 -11372
rect 308 -11520 412 -11321
rect 792 -11372 808 -10948
rect 872 -11372 888 -10948
rect 792 -11388 888 -11372
<< properties >>
string FIXED_BBOX 120 10920 600 11400
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 2 ny 32 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 1 ccov 100
<< end >>
