magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 67 814 203
rect 1 21 697 67
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 177
rect 161 47 191 177
rect 287 47 317 177
rect 383 47 413 177
rect 479 47 509 177
rect 585 47 615 177
rect 696 93 726 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 289 297 325 497
rect 389 297 425 497
rect 483 297 519 497
rect 577 297 613 497
rect 688 297 724 381
<< ndiff >>
rect 27 161 89 177
rect 27 127 35 161
rect 69 127 89 161
rect 27 93 89 127
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 47 161 177
rect 191 89 287 177
rect 191 55 227 89
rect 261 55 287 89
rect 191 47 287 55
rect 317 149 383 177
rect 317 115 337 149
rect 371 115 383 149
rect 317 47 383 115
rect 413 89 479 177
rect 413 55 433 89
rect 467 55 479 89
rect 413 47 479 55
rect 509 165 585 177
rect 509 131 530 165
rect 564 131 585 165
rect 509 47 585 131
rect 615 93 696 177
rect 726 153 788 177
rect 726 119 745 153
rect 779 119 788 153
rect 726 93 788 119
rect 615 89 671 93
rect 615 55 625 89
rect 659 55 671 89
rect 615 47 671 55
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 297 81 451
rect 117 349 175 497
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 489 289 497
rect 211 455 234 489
rect 268 455 289 489
rect 211 297 289 455
rect 325 341 389 497
rect 325 307 343 341
rect 377 307 389 341
rect 325 297 389 307
rect 425 489 483 497
rect 425 455 437 489
rect 471 455 483 489
rect 425 297 483 455
rect 519 341 577 497
rect 519 307 531 341
rect 565 307 577 341
rect 519 297 577 307
rect 613 489 671 497
rect 613 455 625 489
rect 659 455 671 489
rect 613 381 671 455
rect 613 297 688 381
rect 724 356 788 381
rect 724 322 746 356
rect 780 322 788 356
rect 724 297 788 322
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 227 55 261 89
rect 337 115 371 149
rect 433 55 467 89
rect 530 131 564 165
rect 745 119 779 153
rect 625 55 659 89
<< pdiffc >>
rect 35 451 69 485
rect 129 315 163 349
rect 234 455 268 489
rect 343 307 377 341
rect 437 455 471 489
rect 531 307 565 341
rect 625 455 659 489
rect 746 322 780 356
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 289 497 325 523
rect 389 497 425 523
rect 483 497 519 523
rect 577 497 613 523
rect 688 381 724 407
rect 81 282 117 297
rect 175 282 211 297
rect 289 282 325 297
rect 389 282 425 297
rect 483 282 519 297
rect 577 282 613 297
rect 688 282 724 297
rect 79 265 119 282
rect 173 265 213 282
rect 287 265 327 282
rect 387 265 427 282
rect 481 265 521 282
rect 575 265 615 282
rect 686 268 726 282
rect 33 249 119 265
rect 33 215 51 249
rect 85 215 119 249
rect 33 199 119 215
rect 89 177 119 199
rect 161 249 225 265
rect 161 215 171 249
rect 205 215 225 249
rect 161 199 225 215
rect 287 249 615 265
rect 287 215 302 249
rect 336 215 380 249
rect 414 215 615 249
rect 287 199 615 215
rect 657 249 726 268
rect 657 215 667 249
rect 701 215 726 249
rect 657 199 726 215
rect 161 177 191 199
rect 287 177 317 199
rect 383 177 413 199
rect 479 177 509 199
rect 585 177 615 199
rect 696 177 726 199
rect 696 67 726 93
rect 89 21 119 47
rect 161 21 191 47
rect 287 21 317 47
rect 383 21 413 47
rect 479 21 509 47
rect 585 21 615 47
<< polycont >>
rect 51 215 85 249
rect 171 215 205 249
rect 302 215 336 249
rect 380 215 414 249
rect 667 215 701 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 485 85 527
rect 18 451 35 485
rect 69 451 85 485
rect 218 489 284 527
rect 218 455 234 489
rect 268 455 284 489
rect 411 489 487 527
rect 411 455 437 489
rect 471 455 487 489
rect 599 489 675 527
rect 599 455 625 489
rect 659 455 675 489
rect 33 383 788 417
rect 33 265 67 383
rect 745 356 788 383
rect 103 315 129 349
rect 163 315 283 349
rect 103 300 283 315
rect 327 341 596 349
rect 327 307 343 341
rect 377 307 531 341
rect 565 307 596 341
rect 249 297 283 300
rect 249 271 284 297
rect 33 249 85 265
rect 33 215 51 249
rect 33 199 85 215
rect 121 249 215 265
rect 121 215 171 249
rect 205 215 215 249
rect 121 199 215 215
rect 249 249 435 271
rect 249 215 302 249
rect 336 215 380 249
rect 414 215 435 249
rect 249 199 435 215
rect 249 161 291 199
rect 489 165 596 307
rect 18 127 35 161
rect 69 127 291 161
rect 18 123 291 127
rect 335 149 530 165
rect 18 93 85 123
rect 335 115 337 149
rect 371 131 530 149
rect 564 131 596 165
rect 371 123 596 131
rect 640 249 709 349
rect 640 215 667 249
rect 701 215 709 249
rect 640 125 709 215
rect 745 322 746 356
rect 780 322 788 356
rect 745 153 788 322
rect 371 115 373 123
rect 335 99 373 115
rect 779 119 788 153
rect 745 99 788 119
rect 18 59 35 93
rect 69 59 85 93
rect 18 51 85 59
rect 211 55 227 89
rect 261 55 277 89
rect 211 17 277 55
rect 407 55 433 89
rect 467 55 483 89
rect 407 17 483 55
rect 599 55 625 89
rect 659 55 675 89
rect 599 17 675 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 121 221 155 255 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 489 153 523 187 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 673 221 707 255 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and2b_4
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 789080
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 783230
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
