magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 771 203
rect 29 -17 63 21
<< scnmos >>
rect 93 47 123 177
rect 177 47 207 177
rect 365 47 395 177
rect 449 47 479 177
rect 663 47 693 177
<< scpmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 305 297 341 497
rect 451 297 487 497
rect 655 297 691 497
<< ndiff >>
rect 27 161 93 177
rect 27 127 35 161
rect 69 127 93 161
rect 27 93 93 127
rect 27 59 35 93
rect 69 59 93 93
rect 27 47 93 59
rect 123 169 177 177
rect 123 135 133 169
rect 167 135 177 169
rect 123 47 177 135
rect 207 165 259 177
rect 207 131 217 165
rect 251 131 259 165
rect 207 47 259 131
rect 313 93 365 177
rect 313 59 321 93
rect 355 59 365 93
rect 313 47 365 59
rect 395 89 449 177
rect 395 55 405 89
rect 439 55 449 89
rect 395 47 449 55
rect 479 127 537 177
rect 479 93 495 127
rect 529 93 537 127
rect 479 47 537 93
rect 593 169 663 177
rect 593 135 605 169
rect 639 135 663 169
rect 593 101 663 135
rect 593 67 605 101
rect 639 67 663 101
rect 593 47 663 67
rect 693 93 745 177
rect 693 59 703 93
rect 737 59 745 93
rect 693 47 745 59
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 409 179 497
rect 121 375 133 409
rect 167 375 179 409
rect 121 341 179 375
rect 121 307 133 341
rect 167 307 179 341
rect 121 297 179 307
rect 215 297 305 497
rect 341 485 451 497
rect 341 451 379 485
rect 413 451 451 485
rect 341 417 451 451
rect 341 383 379 417
rect 413 383 451 417
rect 341 297 451 383
rect 487 481 541 497
rect 487 447 499 481
rect 533 447 541 481
rect 487 413 541 447
rect 487 379 499 413
rect 533 379 541 413
rect 487 345 541 379
rect 487 311 499 345
rect 533 311 541 345
rect 487 297 541 311
rect 595 477 655 497
rect 595 443 605 477
rect 639 443 655 477
rect 595 409 655 443
rect 595 375 605 409
rect 639 375 655 409
rect 595 297 655 375
rect 691 485 745 497
rect 691 451 703 485
rect 737 451 745 485
rect 691 417 745 451
rect 691 383 703 417
rect 737 383 745 417
rect 691 297 745 383
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 133 135 167 169
rect 217 131 251 165
rect 321 59 355 93
rect 405 55 439 89
rect 495 93 529 127
rect 605 135 639 169
rect 605 67 639 101
rect 703 59 737 93
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 375 167 409
rect 133 307 167 341
rect 379 451 413 485
rect 379 383 413 417
rect 499 447 533 481
rect 499 379 533 413
rect 499 311 533 345
rect 605 443 639 477
rect 605 375 639 409
rect 703 451 737 485
rect 703 383 737 417
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 305 497 341 523
rect 451 497 487 523
rect 655 497 691 523
rect 85 282 121 297
rect 179 282 215 297
rect 305 282 341 297
rect 451 282 487 297
rect 655 282 691 297
rect 83 265 123 282
rect 21 249 123 265
rect 21 215 34 249
rect 68 215 123 249
rect 21 199 123 215
rect 93 177 123 199
rect 177 265 217 282
rect 177 249 248 265
rect 177 215 201 249
rect 235 215 248 249
rect 177 199 248 215
rect 303 259 343 282
rect 449 270 489 282
rect 653 270 693 282
rect 449 265 693 270
rect 303 249 395 259
rect 303 215 319 249
rect 353 215 395 249
rect 303 205 395 215
rect 177 177 207 199
rect 365 177 395 205
rect 449 249 746 265
rect 449 233 701 249
rect 449 177 479 233
rect 663 215 701 233
rect 735 215 746 249
rect 663 198 746 215
rect 663 177 693 198
rect 93 21 123 47
rect 177 21 207 47
rect 365 21 395 47
rect 449 21 479 47
rect 663 21 693 47
<< polycont >>
rect 34 215 68 249
rect 201 215 235 249
rect 319 215 353 249
rect 701 215 735 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 24 477 345 493
rect 24 443 39 477
rect 73 459 345 477
rect 73 443 84 459
rect 24 409 84 443
rect 24 375 39 409
rect 73 375 84 409
rect 24 341 84 375
rect 24 307 39 341
rect 73 307 84 341
rect 24 291 84 307
rect 121 409 178 425
rect 121 375 133 409
rect 167 375 178 409
rect 121 341 178 375
rect 121 307 133 341
rect 167 307 178 341
rect 121 291 178 307
rect 17 249 84 257
rect 17 215 34 249
rect 68 215 84 249
rect 17 212 84 215
rect 17 161 69 177
rect 17 127 35 161
rect 17 93 69 127
rect 121 169 167 291
rect 213 265 253 422
rect 301 330 345 459
rect 379 485 435 527
rect 413 451 435 485
rect 379 417 435 451
rect 413 383 435 417
rect 379 367 435 383
rect 473 481 549 493
rect 473 447 499 481
rect 533 447 549 481
rect 473 413 549 447
rect 473 379 499 413
rect 533 379 549 413
rect 473 345 549 379
rect 473 330 499 345
rect 301 311 499 330
rect 533 311 549 345
rect 301 296 549 311
rect 594 477 639 493
rect 594 443 605 477
rect 594 409 639 443
rect 594 375 605 409
rect 201 249 253 265
rect 594 262 639 375
rect 695 485 754 527
rect 695 451 703 485
rect 737 451 754 485
rect 695 417 754 451
rect 695 383 703 417
rect 737 383 754 417
rect 695 367 754 383
rect 235 215 253 249
rect 297 249 639 262
rect 297 215 319 249
rect 353 215 639 249
rect 201 199 253 215
rect 121 135 133 169
rect 315 165 540 177
rect 121 119 167 135
rect 201 131 217 165
rect 251 143 540 165
rect 251 131 350 143
rect 493 127 540 143
rect 17 59 35 93
rect 69 85 88 93
rect 213 85 321 93
rect 69 59 321 85
rect 355 59 371 93
rect 17 51 371 59
rect 405 89 439 105
rect 405 17 439 55
rect 493 93 495 127
rect 529 93 540 127
rect 493 51 540 93
rect 586 169 639 215
rect 586 135 605 169
rect 673 249 750 324
rect 673 215 701 249
rect 735 215 750 249
rect 673 152 750 215
rect 586 101 639 135
rect 586 67 605 101
rect 586 51 639 67
rect 703 93 747 109
rect 737 59 747 93
rect 703 17 747 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 219 357 253 391 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 703 221 737 255 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 703 153 737 187 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 703 289 737 323 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel locali s 219 289 253 323 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 131 357 165 391 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2i_1
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 1454292
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1447316
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
