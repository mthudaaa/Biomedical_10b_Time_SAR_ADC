magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 8 157 303 203
rect 697 157 897 203
rect 8 67 897 157
rect 29 -17 63 67
rect 305 21 897 67
<< scnmos >>
rect 96 93 126 177
rect 186 93 216 177
rect 393 47 423 131
rect 490 47 520 131
rect 581 47 611 131
rect 678 47 708 131
rect 786 47 816 177
<< scpmoshvt >>
rect 81 410 117 494
rect 385 413 421 497
rect 188 297 224 381
rect 491 297 527 381
rect 573 297 609 381
rect 670 297 706 381
rect 778 297 814 497
<< ndiff >>
rect 34 149 96 177
rect 34 115 42 149
rect 76 115 96 149
rect 34 93 96 115
rect 126 149 186 177
rect 126 115 141 149
rect 175 115 186 149
rect 126 93 186 115
rect 216 149 277 177
rect 216 115 235 149
rect 269 115 277 149
rect 723 131 786 177
rect 216 93 277 115
rect 331 97 393 131
rect 331 63 339 97
rect 373 63 393 97
rect 331 47 393 63
rect 423 111 490 131
rect 423 77 433 111
rect 467 77 490 111
rect 423 47 490 77
rect 520 97 581 131
rect 520 63 530 97
rect 564 63 581 97
rect 520 47 581 63
rect 611 111 678 131
rect 611 77 624 111
rect 658 77 678 111
rect 611 47 678 77
rect 708 97 786 131
rect 708 63 728 97
rect 762 63 786 97
rect 708 47 786 63
rect 816 135 871 177
rect 816 101 826 135
rect 860 101 871 135
rect 816 47 871 101
<< pdiff >>
rect 27 475 81 494
rect 27 441 35 475
rect 69 441 81 475
rect 27 410 81 441
rect 117 475 171 494
rect 117 441 129 475
rect 163 441 171 475
rect 117 410 171 441
rect 331 475 385 497
rect 331 441 339 475
rect 373 441 385 475
rect 331 413 385 441
rect 421 413 474 497
rect 134 381 171 410
rect 134 297 188 381
rect 224 339 282 381
rect 224 305 236 339
rect 270 305 282 339
rect 224 297 282 305
rect 438 381 474 413
rect 723 485 778 497
rect 723 451 731 485
rect 765 451 778 485
rect 723 417 778 451
rect 723 383 731 417
rect 765 383 778 417
rect 723 381 778 383
rect 438 297 491 381
rect 527 297 573 381
rect 609 297 670 381
rect 706 297 778 381
rect 814 454 871 497
rect 814 420 826 454
rect 860 420 871 454
rect 814 386 871 420
rect 814 352 826 386
rect 860 352 871 386
rect 814 297 871 352
<< ndiffc >>
rect 42 115 76 149
rect 141 115 175 149
rect 235 115 269 149
rect 339 63 373 97
rect 433 77 467 111
rect 530 63 564 97
rect 624 77 658 111
rect 728 63 762 97
rect 826 101 860 135
<< pdiffc >>
rect 35 441 69 475
rect 129 441 163 475
rect 339 441 373 475
rect 236 305 270 339
rect 731 451 765 485
rect 731 383 765 417
rect 826 420 860 454
rect 826 352 860 386
<< poly >>
rect 81 494 117 520
rect 385 497 421 523
rect 81 395 117 410
rect 79 265 119 395
rect 188 381 224 407
rect 385 398 421 413
rect 188 282 224 297
rect 186 265 226 282
rect 383 265 423 398
rect 571 484 625 500
rect 778 497 814 523
rect 571 450 581 484
rect 615 450 625 484
rect 571 434 625 450
rect 571 407 611 434
rect 491 381 527 407
rect 573 381 609 407
rect 670 381 706 407
rect 491 282 527 297
rect 573 282 609 297
rect 670 282 706 297
rect 778 282 814 297
rect 489 265 529 282
rect 79 249 133 265
rect 79 215 89 249
rect 123 215 133 249
rect 79 199 133 215
rect 186 249 240 265
rect 186 215 196 249
rect 230 215 240 249
rect 186 199 240 215
rect 367 249 423 265
rect 367 215 377 249
rect 411 215 423 249
rect 367 199 423 215
rect 465 249 529 265
rect 465 215 475 249
rect 509 215 529 249
rect 465 199 529 215
rect 96 177 126 199
rect 186 177 216 199
rect 393 131 423 199
rect 490 131 520 199
rect 571 152 611 282
rect 668 265 708 282
rect 776 265 816 282
rect 654 249 708 265
rect 654 215 664 249
rect 698 215 708 249
rect 654 199 708 215
rect 762 249 816 265
rect 762 215 772 249
rect 806 215 816 249
rect 762 199 816 215
rect 581 131 611 152
rect 678 131 708 199
rect 786 177 816 199
rect 96 67 126 93
rect 186 67 216 93
rect 393 21 423 47
rect 490 21 520 47
rect 581 21 611 47
rect 678 21 708 47
rect 786 21 816 47
<< polycont >>
rect 581 450 615 484
rect 89 215 123 249
rect 196 215 230 249
rect 377 215 411 249
rect 475 215 509 249
rect 664 215 698 249
rect 772 215 806 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 475 69 491
rect 17 441 35 475
rect 103 475 179 527
rect 536 484 674 491
rect 103 441 129 475
rect 163 441 179 475
rect 322 441 339 475
rect 373 441 481 475
rect 17 407 69 441
rect 17 373 403 407
rect 17 165 51 373
rect 85 249 162 339
rect 208 305 236 339
rect 270 305 335 339
rect 85 215 89 249
rect 123 215 162 249
rect 85 199 162 215
rect 196 249 267 265
rect 230 215 267 249
rect 196 199 267 215
rect 301 249 335 305
rect 369 317 403 373
rect 447 391 481 441
rect 536 450 581 484
rect 615 450 674 484
rect 536 425 674 450
rect 718 485 774 527
rect 718 451 731 485
rect 765 451 774 485
rect 718 417 774 451
rect 447 357 674 391
rect 718 383 731 417
rect 765 383 774 417
rect 718 367 774 383
rect 826 454 891 493
rect 860 420 891 454
rect 826 386 891 420
rect 640 333 674 357
rect 860 352 891 386
rect 369 283 509 317
rect 640 299 782 333
rect 826 299 891 352
rect 475 249 509 283
rect 748 265 782 299
rect 301 215 377 249
rect 411 215 431 249
rect 301 165 335 215
rect 475 199 509 215
rect 563 249 714 265
rect 563 215 664 249
rect 698 215 714 249
rect 563 199 714 215
rect 748 249 806 265
rect 748 215 772 249
rect 748 199 806 215
rect 748 165 782 199
rect 17 149 80 165
rect 17 115 42 149
rect 76 115 80 149
rect 17 90 80 115
rect 141 149 175 165
rect 141 17 175 115
rect 235 149 335 165
rect 269 131 335 149
rect 433 131 782 165
rect 847 152 891 299
rect 826 135 891 152
rect 235 90 269 115
rect 433 111 467 131
rect 314 63 339 97
rect 373 63 389 97
rect 314 17 389 63
rect 624 111 658 131
rect 433 61 467 77
rect 504 63 530 97
rect 564 63 580 97
rect 504 17 580 63
rect 860 101 891 135
rect 624 61 658 77
rect 692 63 728 97
rect 762 63 778 97
rect 826 83 891 101
rect 692 17 778 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 563 199 714 265 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 835 357 869 391 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 536 425 674 491 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 196 199 267 265 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 110 221 144 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 or4bb_1
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 2334766
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 2327446
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
