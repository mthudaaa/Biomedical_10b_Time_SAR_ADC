magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 1 67 1282 203
rect 29 -17 63 67
rect 301 21 1282 67
<< scnmos >>
rect 79 93 109 177
rect 186 93 216 177
rect 405 47 435 177
rect 499 47 529 177
rect 583 47 613 177
rect 687 47 717 177
rect 879 47 909 177
rect 983 47 1013 177
rect 1067 47 1097 177
rect 1171 47 1201 177
<< scpmoshvt >>
rect 81 410 117 494
rect 188 297 224 381
rect 397 297 433 497
rect 491 297 527 497
rect 585 297 621 497
rect 679 297 715 497
rect 881 297 917 497
rect 975 297 1011 497
rect 1069 297 1105 497
rect 1163 297 1199 497
<< ndiff >>
rect 27 149 79 177
rect 27 115 35 149
rect 69 115 79 149
rect 27 93 79 115
rect 109 149 186 177
rect 109 115 137 149
rect 171 115 186 149
rect 109 93 186 115
rect 216 149 273 177
rect 216 115 231 149
rect 265 115 273 149
rect 216 93 273 115
rect 327 95 405 177
rect 327 61 335 95
rect 369 61 405 95
rect 327 47 405 61
rect 435 163 499 177
rect 435 129 445 163
rect 479 129 499 163
rect 435 95 499 129
rect 435 61 445 95
rect 479 61 499 95
rect 435 47 499 61
rect 529 95 583 177
rect 529 61 539 95
rect 573 61 583 95
rect 529 47 583 61
rect 613 163 687 177
rect 613 129 633 163
rect 667 129 687 163
rect 613 95 687 129
rect 613 61 633 95
rect 667 61 687 95
rect 613 47 687 61
rect 717 95 769 177
rect 717 61 727 95
rect 761 61 769 95
rect 717 47 769 61
rect 823 95 879 177
rect 823 61 835 95
rect 869 61 879 95
rect 823 47 879 61
rect 909 163 983 177
rect 909 129 929 163
rect 963 129 983 163
rect 909 95 983 129
rect 909 61 929 95
rect 963 61 983 95
rect 909 47 983 61
rect 1013 95 1067 177
rect 1013 61 1023 95
rect 1057 61 1067 95
rect 1013 47 1067 61
rect 1097 163 1171 177
rect 1097 129 1117 163
rect 1151 129 1171 163
rect 1097 95 1171 129
rect 1097 61 1117 95
rect 1151 61 1171 95
rect 1097 47 1171 61
rect 1201 163 1256 177
rect 1201 129 1211 163
rect 1245 129 1256 163
rect 1201 95 1256 129
rect 1201 61 1211 95
rect 1245 61 1256 95
rect 1201 47 1256 61
<< pdiff >>
rect 27 475 81 494
rect 27 441 35 475
rect 69 441 81 475
rect 27 410 81 441
rect 117 482 171 494
rect 117 448 129 482
rect 163 448 171 482
rect 117 410 171 448
rect 134 381 171 410
rect 343 479 397 497
rect 343 445 351 479
rect 385 445 397 479
rect 134 297 188 381
rect 224 343 278 381
rect 224 309 236 343
rect 270 309 278 343
rect 224 297 278 309
rect 343 297 397 445
rect 433 409 491 497
rect 433 375 445 409
rect 479 375 491 409
rect 433 297 491 375
rect 527 479 585 497
rect 527 445 539 479
rect 573 445 585 479
rect 527 297 585 445
rect 621 341 679 497
rect 621 307 633 341
rect 667 307 679 341
rect 621 297 679 307
rect 715 479 769 497
rect 715 445 727 479
rect 761 445 769 479
rect 715 297 769 445
rect 823 477 881 497
rect 823 443 835 477
rect 869 443 881 477
rect 823 297 881 443
rect 917 409 975 497
rect 917 375 929 409
rect 963 375 975 409
rect 917 341 975 375
rect 917 307 929 341
rect 963 307 975 341
rect 917 297 975 307
rect 1011 477 1069 497
rect 1011 443 1023 477
rect 1057 443 1069 477
rect 1011 409 1069 443
rect 1011 375 1023 409
rect 1057 375 1069 409
rect 1011 341 1069 375
rect 1011 307 1023 341
rect 1057 307 1069 341
rect 1011 297 1069 307
rect 1105 477 1163 497
rect 1105 443 1117 477
rect 1151 443 1163 477
rect 1105 409 1163 443
rect 1105 375 1117 409
rect 1151 375 1163 409
rect 1105 297 1163 375
rect 1199 479 1256 497
rect 1199 445 1211 479
rect 1245 445 1256 479
rect 1199 411 1256 445
rect 1199 377 1211 411
rect 1245 377 1256 411
rect 1199 343 1256 377
rect 1199 309 1211 343
rect 1245 309 1256 343
rect 1199 297 1256 309
<< ndiffc >>
rect 35 115 69 149
rect 137 115 171 149
rect 231 115 265 149
rect 335 61 369 95
rect 445 129 479 163
rect 445 61 479 95
rect 539 61 573 95
rect 633 129 667 163
rect 633 61 667 95
rect 727 61 761 95
rect 835 61 869 95
rect 929 129 963 163
rect 929 61 963 95
rect 1023 61 1057 95
rect 1117 129 1151 163
rect 1117 61 1151 95
rect 1211 129 1245 163
rect 1211 61 1245 95
<< pdiffc >>
rect 35 441 69 475
rect 129 448 163 482
rect 351 445 385 479
rect 236 309 270 343
rect 445 375 479 409
rect 539 445 573 479
rect 633 307 667 341
rect 727 445 761 479
rect 835 443 869 477
rect 929 375 963 409
rect 929 307 963 341
rect 1023 443 1057 477
rect 1023 375 1057 409
rect 1023 307 1057 341
rect 1117 443 1151 477
rect 1117 375 1151 409
rect 1211 445 1245 479
rect 1211 377 1245 411
rect 1211 309 1245 343
<< poly >>
rect 81 494 117 520
rect 397 497 433 523
rect 491 497 527 523
rect 585 497 621 523
rect 679 497 715 523
rect 881 497 917 523
rect 975 497 1011 523
rect 1069 497 1105 523
rect 1163 497 1199 523
rect 81 395 117 410
rect 79 265 119 395
rect 188 381 224 407
rect 188 282 224 297
rect 397 282 433 297
rect 491 282 527 297
rect 585 282 621 297
rect 679 282 715 297
rect 881 282 917 297
rect 975 282 1011 297
rect 1069 282 1105 297
rect 1163 282 1199 297
rect 186 265 226 282
rect 395 265 435 282
rect 489 265 529 282
rect 79 249 139 265
rect 79 215 89 249
rect 123 215 139 249
rect 79 199 139 215
rect 186 249 260 265
rect 186 215 200 249
rect 234 215 260 249
rect 186 199 260 215
rect 357 249 529 265
rect 357 215 367 249
rect 401 215 445 249
rect 479 215 529 249
rect 357 199 529 215
rect 79 177 109 199
rect 186 177 216 199
rect 405 177 435 199
rect 499 177 529 199
rect 583 265 623 282
rect 677 265 717 282
rect 583 249 717 265
rect 583 215 593 249
rect 627 215 671 249
rect 705 215 717 249
rect 583 199 717 215
rect 583 177 613 199
rect 687 177 717 199
rect 879 265 919 282
rect 973 265 1013 282
rect 879 249 1013 265
rect 879 215 932 249
rect 966 215 1013 249
rect 879 199 1013 215
rect 879 177 909 199
rect 983 177 1013 199
rect 1067 265 1107 282
rect 1161 265 1201 282
rect 1067 249 1201 265
rect 1067 215 1119 249
rect 1153 215 1201 249
rect 1067 199 1201 215
rect 1067 177 1097 199
rect 1171 177 1201 199
rect 79 67 109 93
rect 186 67 216 93
rect 405 21 435 47
rect 499 21 529 47
rect 583 21 613 47
rect 687 21 717 47
rect 879 21 909 47
rect 983 21 1013 47
rect 1067 21 1097 47
rect 1171 21 1201 47
<< polycont >>
rect 89 215 123 249
rect 200 215 234 249
rect 367 215 401 249
rect 445 215 479 249
rect 593 215 627 249
rect 671 215 705 249
rect 932 215 966 249
rect 1119 215 1153 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 475 69 491
rect 17 441 35 475
rect 103 482 179 527
rect 103 448 129 482
rect 163 448 179 482
rect 335 479 777 493
rect 335 445 351 479
rect 385 445 539 479
rect 573 445 727 479
rect 761 445 777 479
rect 819 477 1065 493
rect 819 443 835 477
rect 869 443 1023 477
rect 1057 443 1065 477
rect 17 411 69 441
rect 17 377 390 411
rect 1023 409 1065 443
rect 17 165 51 377
rect 85 249 166 339
rect 209 309 236 343
rect 270 309 322 343
rect 209 305 322 309
rect 85 215 89 249
rect 123 215 166 249
rect 85 199 166 215
rect 200 249 254 265
rect 234 215 254 249
rect 200 199 254 215
rect 288 249 322 305
rect 356 317 390 377
rect 429 375 445 409
rect 479 375 929 409
rect 963 375 979 409
rect 921 341 979 375
rect 356 283 573 317
rect 607 307 633 341
rect 667 307 846 341
rect 607 289 846 307
rect 921 307 929 341
rect 963 307 979 341
rect 921 291 979 307
rect 1057 375 1065 409
rect 1023 341 1065 375
rect 1109 477 1151 527
rect 1109 443 1117 477
rect 1109 409 1151 443
rect 1109 375 1117 409
rect 1109 359 1151 375
rect 1185 479 1261 493
rect 1185 445 1211 479
rect 1245 445 1261 479
rect 1185 411 1261 445
rect 1185 377 1211 411
rect 1245 377 1261 411
rect 1057 325 1065 341
rect 1185 343 1261 377
rect 1185 325 1211 343
rect 1057 309 1211 325
rect 1245 309 1261 343
rect 1057 307 1261 309
rect 1023 291 1261 307
rect 539 255 573 283
rect 539 249 728 255
rect 288 215 367 249
rect 401 215 445 249
rect 479 215 495 249
rect 539 215 593 249
rect 627 215 671 249
rect 705 215 728 249
rect 288 165 322 215
rect 762 181 846 289
rect 880 249 1059 255
rect 880 215 932 249
rect 966 215 1059 249
rect 1093 249 1266 255
rect 1093 215 1119 249
rect 1153 215 1266 249
rect 17 149 93 165
rect 17 115 35 149
rect 69 115 93 149
rect 17 90 93 115
rect 137 149 171 165
rect 137 17 171 115
rect 231 149 322 165
rect 265 131 322 149
rect 419 163 1167 181
rect 265 115 270 131
rect 231 90 270 115
rect 419 129 445 163
rect 479 145 633 163
rect 479 129 495 145
rect 319 95 385 96
rect 319 61 335 95
rect 369 61 385 95
rect 319 17 385 61
rect 419 95 495 129
rect 607 129 633 145
rect 667 145 929 163
rect 667 129 683 145
rect 419 61 445 95
rect 479 61 495 95
rect 419 51 495 61
rect 539 95 573 111
rect 539 17 573 61
rect 607 95 683 129
rect 903 129 929 145
rect 963 145 1117 163
rect 963 129 979 145
rect 607 61 633 95
rect 667 61 683 95
rect 607 51 683 61
rect 727 95 869 111
rect 761 61 835 95
rect 727 17 869 61
rect 903 95 979 129
rect 1091 129 1117 145
rect 1151 129 1167 163
rect 903 61 929 95
rect 963 61 979 95
rect 903 51 979 61
rect 1023 95 1057 111
rect 1023 17 1057 61
rect 1091 95 1167 129
rect 1091 61 1117 95
rect 1151 61 1167 95
rect 1091 51 1167 61
rect 1211 163 1266 181
rect 1245 129 1266 163
rect 1211 95 1266 129
rect 1245 61 1266 95
rect 1211 17 1266 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 132 221 166 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 210 221 244 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel locali s 1118 221 1152 255 0 FreeSans 400 180 0 0 A
port 1 nsew signal input
flabel locali s 720 289 754 323 0 FreeSans 400 180 0 0 Y
port 9 nsew signal output
flabel locali s 914 221 948 255 0 FreeSans 400 180 0 0 B
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 -10 0 -10 4 nor4bb_2
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 1835486
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1825954
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
