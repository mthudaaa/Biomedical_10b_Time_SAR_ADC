magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 725 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 174 47 204 177
rect 384 47 414 177
rect 470 47 500 177
rect 606 47 636 177
<< scpmoshvt >>
rect 81 297 117 497
rect 176 297 212 497
rect 376 297 412 497
rect 472 297 508 497
rect 608 297 644 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 101 174 177
rect 109 67 129 101
rect 163 67 174 101
rect 109 47 174 67
rect 204 93 267 177
rect 204 59 225 93
rect 259 59 267 93
rect 204 47 267 59
rect 321 162 384 177
rect 321 128 329 162
rect 363 128 384 162
rect 321 94 384 128
rect 321 60 329 94
rect 363 60 384 94
rect 321 47 384 60
rect 414 149 470 177
rect 414 115 425 149
rect 459 115 470 149
rect 414 47 470 115
rect 500 93 606 177
rect 500 59 525 93
rect 559 59 606 93
rect 500 47 606 59
rect 636 149 699 177
rect 636 115 657 149
rect 691 115 699 149
rect 636 47 699 115
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 380 81 451
rect 27 346 35 380
rect 69 346 81 380
rect 27 297 81 346
rect 117 477 176 497
rect 117 443 129 477
rect 163 443 176 477
rect 117 379 176 443
rect 117 345 129 379
rect 163 345 176 379
rect 117 297 176 345
rect 212 485 376 497
rect 212 451 225 485
rect 259 451 329 485
rect 363 451 376 485
rect 212 297 376 451
rect 412 477 472 497
rect 412 443 425 477
rect 459 443 472 477
rect 412 401 472 443
rect 412 367 425 401
rect 459 367 472 401
rect 412 297 472 367
rect 508 297 608 497
rect 644 485 699 497
rect 644 451 657 485
rect 691 451 699 485
rect 644 385 699 451
rect 644 351 657 385
rect 691 351 699 385
rect 644 297 699 351
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 67 163 101
rect 225 59 259 93
rect 329 128 363 162
rect 329 60 363 94
rect 425 115 459 149
rect 525 59 559 93
rect 657 115 691 149
<< pdiffc >>
rect 35 451 69 485
rect 35 346 69 380
rect 129 443 163 477
rect 129 345 163 379
rect 225 451 259 485
rect 329 451 363 485
rect 425 443 459 477
rect 425 367 459 401
rect 657 451 691 485
rect 657 351 691 385
<< poly >>
rect 81 497 117 523
rect 176 497 212 523
rect 376 497 412 523
rect 472 497 508 523
rect 608 497 644 523
rect 81 282 117 297
rect 176 282 212 297
rect 376 282 412 297
rect 472 282 508 297
rect 608 282 644 297
rect 79 267 119 282
rect 174 267 214 282
rect 79 265 214 267
rect 374 265 414 282
rect 79 249 243 265
rect 79 215 199 249
rect 233 215 243 249
rect 79 199 243 215
rect 325 249 414 265
rect 325 215 341 249
rect 375 215 414 249
rect 325 199 414 215
rect 79 177 109 199
rect 174 177 204 199
rect 384 177 414 199
rect 470 265 510 282
rect 606 265 646 282
rect 470 249 532 265
rect 470 215 480 249
rect 514 215 532 249
rect 470 199 532 215
rect 606 249 704 265
rect 606 215 660 249
rect 694 215 704 249
rect 606 199 704 215
rect 470 177 500 199
rect 606 177 636 199
rect 79 21 109 47
rect 174 21 204 47
rect 384 21 414 47
rect 470 21 500 47
rect 606 21 636 47
<< polycont >>
rect 199 215 233 249
rect 341 215 375 249
rect 480 215 514 249
rect 660 215 694 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 380 69 451
rect 18 346 35 380
rect 18 327 69 346
rect 106 477 165 493
rect 106 443 129 477
rect 163 443 165 477
rect 106 379 165 443
rect 199 485 379 527
rect 199 451 225 485
rect 259 451 329 485
rect 363 451 379 485
rect 199 437 379 451
rect 423 477 475 493
rect 423 443 425 477
rect 459 443 475 477
rect 423 401 475 443
rect 106 345 129 379
rect 163 345 165 379
rect 21 161 69 177
rect 21 127 35 161
rect 21 93 69 127
rect 21 59 35 93
rect 21 17 69 59
rect 106 101 165 345
rect 237 367 425 401
rect 459 367 475 401
rect 649 485 706 527
rect 649 451 657 485
rect 691 451 706 485
rect 237 357 475 367
rect 237 266 271 357
rect 199 249 271 266
rect 233 215 271 249
rect 199 168 271 215
rect 305 249 391 323
rect 560 280 615 397
rect 649 385 706 451
rect 649 351 657 385
rect 691 351 706 385
rect 649 330 706 351
rect 305 215 341 249
rect 375 215 391 249
rect 305 202 391 215
rect 464 249 615 280
rect 464 215 480 249
rect 514 215 615 249
rect 464 205 615 215
rect 655 249 707 290
rect 655 215 660 249
rect 694 215 707 249
rect 655 199 707 215
rect 199 162 379 168
rect 199 128 329 162
rect 363 128 379 162
rect 199 127 379 128
rect 106 67 129 101
rect 163 67 165 101
rect 313 94 379 127
rect 106 51 165 67
rect 199 59 225 93
rect 259 59 275 93
rect 199 17 275 59
rect 313 60 329 94
rect 363 60 379 94
rect 423 149 706 165
rect 423 115 425 149
rect 459 127 657 149
rect 459 115 465 127
rect 423 93 465 115
rect 651 115 657 127
rect 691 115 706 149
rect 651 99 706 115
rect 313 51 379 60
rect 499 59 525 93
rect 559 59 607 93
rect 499 17 607 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 662 221 696 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 305 202 391 323 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 580 357 614 391 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 130 425 164 459 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21a_2
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 1908980
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1903184
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
