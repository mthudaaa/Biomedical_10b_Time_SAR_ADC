magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -65 261 1234 582
<< pwell >>
rect 1 21 1151 203
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 177
rect 173 47 203 177
rect 277 47 307 177
rect 371 47 401 177
rect 455 47 485 177
rect 549 47 579 177
rect 747 47 777 177
rect 851 47 881 177
rect 935 47 965 177
rect 1039 47 1069 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 749 297 785 497
rect 843 297 879 497
rect 937 297 973 497
rect 1031 297 1067 497
<< ndiff >>
rect 27 163 89 177
rect 27 129 35 163
rect 69 129 89 163
rect 27 95 89 129
rect 27 61 35 95
rect 69 61 89 95
rect 27 47 89 61
rect 119 163 173 177
rect 119 129 129 163
rect 163 129 173 163
rect 119 95 173 129
rect 119 61 129 95
rect 163 61 173 95
rect 119 47 173 61
rect 203 163 277 177
rect 203 129 223 163
rect 257 129 277 163
rect 203 47 277 129
rect 307 95 371 177
rect 307 61 317 95
rect 351 61 371 95
rect 307 47 371 61
rect 401 95 455 177
rect 401 61 411 95
rect 445 61 455 95
rect 401 47 455 61
rect 485 163 549 177
rect 485 129 505 163
rect 539 129 549 163
rect 485 95 549 129
rect 485 61 505 95
rect 539 61 549 95
rect 485 47 549 61
rect 579 95 747 177
rect 579 61 599 95
rect 633 61 703 95
rect 737 61 747 95
rect 579 47 747 61
rect 777 163 851 177
rect 777 129 797 163
rect 831 129 851 163
rect 777 95 851 129
rect 777 61 797 95
rect 831 61 851 95
rect 777 47 851 61
rect 881 95 935 177
rect 881 61 891 95
rect 925 61 935 95
rect 881 47 935 61
rect 965 163 1039 177
rect 965 129 985 163
rect 1019 129 1039 163
rect 965 95 1039 129
rect 965 61 985 95
rect 1019 61 1039 95
rect 965 47 1039 61
rect 1069 163 1125 177
rect 1069 129 1079 163
rect 1113 129 1125 163
rect 1069 95 1125 129
rect 1069 61 1079 95
rect 1113 61 1125 95
rect 1069 47 1125 61
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 297 81 375
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 297 175 443
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 409 269 443
rect 211 375 223 409
rect 257 375 269 409
rect 211 297 269 375
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 297 363 443
rect 399 477 457 497
rect 399 443 411 477
rect 445 443 457 477
rect 399 409 457 443
rect 399 375 411 409
rect 445 375 457 409
rect 399 297 457 375
rect 493 409 551 497
rect 493 375 505 409
rect 539 375 551 409
rect 493 341 551 375
rect 493 307 505 341
rect 539 307 551 341
rect 493 297 551 307
rect 587 477 641 497
rect 587 443 599 477
rect 633 443 641 477
rect 587 409 641 443
rect 587 375 599 409
rect 633 375 641 409
rect 587 297 641 375
rect 695 477 749 497
rect 695 443 703 477
rect 737 443 749 477
rect 695 409 749 443
rect 695 375 703 409
rect 737 375 749 409
rect 695 297 749 375
rect 785 477 843 497
rect 785 443 797 477
rect 831 443 843 477
rect 785 297 843 443
rect 879 477 937 497
rect 879 443 891 477
rect 925 443 937 477
rect 879 409 937 443
rect 879 375 891 409
rect 925 375 937 409
rect 879 297 937 375
rect 973 409 1031 497
rect 973 375 985 409
rect 1019 375 1031 409
rect 973 341 1031 375
rect 973 307 985 341
rect 1019 307 1031 341
rect 973 297 1031 307
rect 1067 477 1125 497
rect 1067 443 1079 477
rect 1113 443 1125 477
rect 1067 409 1125 443
rect 1067 375 1079 409
rect 1113 375 1125 409
rect 1067 341 1125 375
rect 1067 307 1079 341
rect 1113 307 1125 341
rect 1067 297 1125 307
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 129 129 163 163
rect 129 61 163 95
rect 223 129 257 163
rect 317 61 351 95
rect 411 61 445 95
rect 505 129 539 163
rect 505 61 539 95
rect 599 61 633 95
rect 703 61 737 95
rect 797 129 831 163
rect 797 61 831 95
rect 891 61 925 95
rect 985 129 1019 163
rect 985 61 1019 95
rect 1079 129 1113 163
rect 1079 61 1113 95
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 443 163 477
rect 223 443 257 477
rect 223 375 257 409
rect 317 443 351 477
rect 411 443 445 477
rect 411 375 445 409
rect 505 375 539 409
rect 505 307 539 341
rect 599 443 633 477
rect 599 375 633 409
rect 703 443 737 477
rect 703 375 737 409
rect 797 443 831 477
rect 891 443 925 477
rect 891 375 925 409
rect 985 375 1019 409
rect 985 307 1019 341
rect 1079 443 1113 477
rect 1079 375 1113 409
rect 1079 307 1113 341
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 749 497 785 523
rect 843 497 879 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 749 282 785 297
rect 843 282 879 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 79 265 119 282
rect 55 249 119 265
rect 55 215 65 249
rect 99 215 119 249
rect 55 199 119 215
rect 89 177 119 199
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 747 265 787 282
rect 841 265 881 282
rect 173 249 307 265
rect 173 215 223 249
rect 257 215 307 249
rect 173 199 307 215
rect 349 249 413 265
rect 349 215 359 249
rect 393 215 413 249
rect 349 199 413 215
rect 455 249 649 265
rect 455 215 599 249
rect 633 215 649 249
rect 455 199 649 215
rect 747 249 881 265
rect 747 215 795 249
rect 829 215 881 249
rect 747 199 881 215
rect 173 177 203 199
rect 277 177 307 199
rect 371 177 401 199
rect 455 177 485 199
rect 549 177 579 199
rect 747 177 777 199
rect 851 177 881 199
rect 935 265 975 282
rect 1029 265 1069 282
rect 935 249 1069 265
rect 935 215 987 249
rect 1021 215 1069 249
rect 935 199 1069 215
rect 935 177 965 199
rect 1039 177 1069 199
rect 89 21 119 47
rect 173 21 203 47
rect 277 21 307 47
rect 371 21 401 47
rect 455 21 485 47
rect 549 21 579 47
rect 747 21 777 47
rect 851 21 881 47
rect 935 21 965 47
rect 1039 21 1069 47
<< polycont >>
rect 65 215 99 249
rect 223 215 257 249
rect 359 215 393 249
rect 599 215 633 249
rect 795 215 829 249
rect 987 215 1021 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 27 477 77 493
rect 27 443 35 477
rect 69 443 77 477
rect 27 409 77 443
rect 121 477 171 527
rect 121 443 129 477
rect 163 443 171 477
rect 121 427 171 443
rect 215 477 265 493
rect 215 443 223 477
rect 257 443 265 477
rect 27 375 35 409
rect 69 391 77 409
rect 215 409 265 443
rect 309 477 359 527
rect 309 443 317 477
rect 351 443 359 477
rect 309 427 359 443
rect 403 477 641 493
rect 403 443 411 477
rect 445 459 599 477
rect 445 443 453 459
rect 215 391 223 409
rect 69 375 223 391
rect 257 391 265 409
rect 403 409 453 443
rect 591 443 599 459
rect 633 443 641 477
rect 403 391 411 409
rect 257 375 411 391
rect 445 375 453 409
rect 27 357 453 375
rect 489 409 555 425
rect 489 375 505 409
rect 539 375 555 409
rect 489 341 555 375
rect 591 409 641 443
rect 591 375 599 409
rect 633 375 641 409
rect 591 359 641 375
rect 695 477 745 493
rect 695 443 703 477
rect 737 443 745 477
rect 695 409 745 443
rect 789 477 839 527
rect 789 443 797 477
rect 831 443 839 477
rect 789 427 839 443
rect 883 477 1121 493
rect 883 443 891 477
rect 925 459 1079 477
rect 925 443 933 459
rect 695 375 703 409
rect 737 393 745 409
rect 883 409 933 443
rect 1071 443 1079 459
rect 1113 443 1121 477
rect 883 393 891 409
rect 737 375 891 393
rect 925 375 933 409
rect 695 357 933 375
rect 977 409 1027 425
rect 977 375 985 409
rect 1019 375 1027 409
rect 22 289 419 323
rect 22 249 128 289
rect 22 215 65 249
rect 99 215 128 249
rect 171 249 289 255
rect 171 215 223 249
rect 257 215 289 249
rect 343 249 419 289
rect 343 215 359 249
rect 393 215 419 249
rect 489 307 505 341
rect 539 307 555 341
rect 977 341 1027 375
rect 977 323 985 341
rect 489 181 555 307
rect 623 307 985 323
rect 1019 307 1027 341
rect 623 289 1027 307
rect 1071 409 1121 443
rect 1071 375 1079 409
rect 1113 375 1121 409
rect 1071 341 1121 375
rect 1071 307 1079 341
rect 1113 307 1121 341
rect 1071 291 1121 307
rect 623 265 657 289
rect 599 249 657 265
rect 633 215 657 249
rect 695 249 894 255
rect 695 215 795 249
rect 829 215 894 249
rect 944 249 1087 255
rect 944 215 987 249
rect 1021 215 1087 249
rect 599 199 657 215
rect 35 163 69 179
rect 35 95 69 129
rect 35 17 69 61
rect 103 163 163 179
rect 103 129 129 163
rect 197 163 555 181
rect 197 129 223 163
rect 257 145 505 163
rect 257 129 273 145
rect 479 129 505 145
rect 539 129 555 163
rect 623 181 657 199
rect 623 163 1035 181
rect 623 145 797 163
rect 103 95 163 129
rect 411 95 445 111
rect 103 61 129 95
rect 163 61 317 95
rect 351 61 367 95
rect 103 51 367 61
rect 411 17 445 61
rect 479 95 555 129
rect 771 129 797 145
rect 831 145 985 163
rect 831 129 847 145
rect 479 61 505 95
rect 539 61 555 95
rect 479 51 555 61
rect 599 95 737 111
rect 633 61 703 95
rect 599 17 737 61
rect 771 95 847 129
rect 959 129 985 145
rect 1019 129 1035 163
rect 771 61 797 95
rect 831 61 847 95
rect 771 51 847 61
rect 891 95 925 111
rect 891 17 925 61
rect 959 95 1035 129
rect 959 61 985 95
rect 1019 61 1035 95
rect 959 51 1035 61
rect 1079 163 1113 181
rect 1079 95 1113 129
rect 1079 17 1113 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 1016 221 1050 255 0 FreeSans 400 180 0 0 A2_N
port 2 nsew signal input
flabel locali s 695 215 894 255 0 FreeSans 400 180 0 0 A1_N
port 1 nsew signal input
flabel locali s 512 289 546 323 0 FreeSans 400 180 0 0 Y
port 9 nsew signal output
flabel locali s 196 221 230 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 62 221 96 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2bb2oi_2
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 523626
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 514428
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
