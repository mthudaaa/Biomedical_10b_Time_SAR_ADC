magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 23 21 1517 203
rect 29 -17 63 21
<< scnmos >>
rect 101 47 131 177
rect 183 47 213 177
rect 267 47 297 177
rect 349 47 379 177
rect 465 47 495 177
rect 549 47 579 177
rect 757 47 787 177
rect 841 47 871 177
rect 945 47 975 177
rect 1029 47 1059 177
rect 1133 47 1163 177
rect 1217 47 1247 177
rect 1321 47 1351 177
rect 1405 47 1435 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 749 297 785 497
rect 843 297 879 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1125 297 1161 497
rect 1219 297 1255 497
rect 1313 297 1349 497
rect 1407 297 1443 497
<< ndiff >>
rect 49 161 101 177
rect 49 127 57 161
rect 91 127 101 161
rect 49 93 101 127
rect 49 59 57 93
rect 91 59 101 93
rect 49 47 101 59
rect 131 47 183 177
rect 213 165 267 177
rect 213 131 223 165
rect 257 131 267 165
rect 213 93 267 131
rect 213 59 223 93
rect 257 59 267 93
rect 213 47 267 59
rect 297 47 349 177
rect 379 93 465 177
rect 379 59 405 93
rect 439 59 465 93
rect 379 47 465 59
rect 495 169 549 177
rect 495 135 505 169
rect 539 135 549 169
rect 495 101 549 135
rect 495 67 505 101
rect 539 67 549 101
rect 495 47 549 67
rect 579 93 757 177
rect 579 59 599 93
rect 633 59 697 93
rect 731 59 757 93
rect 579 47 757 59
rect 787 165 841 177
rect 787 131 797 165
rect 831 131 841 165
rect 787 89 841 131
rect 787 55 797 89
rect 831 55 841 89
rect 787 47 841 55
rect 871 89 945 177
rect 871 55 891 89
rect 925 55 945 89
rect 871 47 945 55
rect 975 165 1029 177
rect 975 131 985 165
rect 1019 131 1029 165
rect 975 89 1029 131
rect 975 55 985 89
rect 1019 55 1029 89
rect 975 47 1029 55
rect 1059 89 1133 177
rect 1059 55 1079 89
rect 1113 55 1133 89
rect 1059 47 1133 55
rect 1163 165 1217 177
rect 1163 131 1173 165
rect 1207 131 1217 165
rect 1163 89 1217 131
rect 1163 55 1173 89
rect 1207 55 1217 89
rect 1163 47 1217 55
rect 1247 89 1321 177
rect 1247 55 1267 89
rect 1301 55 1321 89
rect 1247 47 1321 55
rect 1351 165 1405 177
rect 1351 131 1361 165
rect 1395 131 1405 165
rect 1351 89 1405 131
rect 1351 55 1361 89
rect 1395 55 1405 89
rect 1351 47 1405 55
rect 1435 165 1491 177
rect 1435 131 1445 165
rect 1479 131 1491 165
rect 1435 89 1491 131
rect 1435 55 1445 89
rect 1479 55 1491 89
rect 1435 47 1491 55
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 478 175 497
rect 117 444 129 478
rect 163 444 175 478
rect 117 297 175 444
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 394 269 443
rect 211 360 223 394
rect 257 360 269 394
rect 211 297 269 360
rect 305 478 363 497
rect 305 444 317 478
rect 351 444 363 478
rect 305 297 363 444
rect 399 479 457 497
rect 399 445 411 479
rect 445 445 457 479
rect 399 411 457 445
rect 399 377 411 411
rect 445 377 457 411
rect 399 343 457 377
rect 399 309 411 343
rect 445 309 457 343
rect 399 297 457 309
rect 493 409 551 497
rect 493 375 505 409
rect 539 375 551 409
rect 493 341 551 375
rect 493 307 505 341
rect 539 307 551 341
rect 493 297 551 307
rect 587 485 641 497
rect 587 451 599 485
rect 633 451 641 485
rect 587 391 641 451
rect 587 357 599 391
rect 633 357 641 391
rect 587 297 641 357
rect 695 485 749 497
rect 695 451 703 485
rect 737 451 749 485
rect 695 417 749 451
rect 695 383 703 417
rect 737 383 749 417
rect 695 349 749 383
rect 695 315 703 349
rect 737 315 749 349
rect 695 297 749 315
rect 785 477 843 497
rect 785 443 797 477
rect 831 443 843 477
rect 785 409 843 443
rect 785 375 797 409
rect 831 375 843 409
rect 785 341 843 375
rect 785 307 797 341
rect 831 307 843 341
rect 785 297 843 307
rect 879 489 937 497
rect 879 455 891 489
rect 925 455 937 489
rect 879 391 937 455
rect 879 357 891 391
rect 925 357 937 391
rect 879 297 937 357
rect 973 477 1031 497
rect 973 443 985 477
rect 1019 443 1031 477
rect 973 409 1031 443
rect 973 375 985 409
rect 1019 375 1031 409
rect 973 341 1031 375
rect 973 307 985 341
rect 1019 307 1031 341
rect 973 297 1031 307
rect 1067 489 1125 497
rect 1067 455 1079 489
rect 1113 455 1125 489
rect 1067 391 1125 455
rect 1067 357 1079 391
rect 1113 357 1125 391
rect 1067 297 1125 357
rect 1161 477 1219 497
rect 1161 443 1173 477
rect 1207 443 1219 477
rect 1161 409 1219 443
rect 1161 375 1173 409
rect 1207 375 1219 409
rect 1161 341 1219 375
rect 1161 307 1173 341
rect 1207 307 1219 341
rect 1161 297 1219 307
rect 1255 489 1313 497
rect 1255 455 1267 489
rect 1301 455 1313 489
rect 1255 391 1313 455
rect 1255 357 1267 391
rect 1301 357 1313 391
rect 1255 297 1313 357
rect 1349 477 1407 497
rect 1349 443 1361 477
rect 1395 443 1407 477
rect 1349 409 1407 443
rect 1349 375 1361 409
rect 1395 375 1407 409
rect 1349 341 1407 375
rect 1349 307 1361 341
rect 1395 307 1407 341
rect 1349 297 1407 307
rect 1443 479 1497 497
rect 1443 445 1455 479
rect 1489 445 1497 479
rect 1443 411 1497 445
rect 1443 377 1455 411
rect 1489 377 1497 411
rect 1443 343 1497 377
rect 1443 309 1455 343
rect 1489 309 1497 343
rect 1443 297 1497 309
<< ndiffc >>
rect 57 127 91 161
rect 57 59 91 93
rect 223 131 257 165
rect 223 59 257 93
rect 405 59 439 93
rect 505 135 539 169
rect 505 67 539 101
rect 599 59 633 93
rect 697 59 731 93
rect 797 131 831 165
rect 797 55 831 89
rect 891 55 925 89
rect 985 131 1019 165
rect 985 55 1019 89
rect 1079 55 1113 89
rect 1173 131 1207 165
rect 1173 55 1207 89
rect 1267 55 1301 89
rect 1361 131 1395 165
rect 1361 55 1395 89
rect 1445 131 1479 165
rect 1445 55 1479 89
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 444 163 478
rect 223 443 257 477
rect 223 360 257 394
rect 317 444 351 478
rect 411 445 445 479
rect 411 377 445 411
rect 411 309 445 343
rect 505 375 539 409
rect 505 307 539 341
rect 599 451 633 485
rect 599 357 633 391
rect 703 451 737 485
rect 703 383 737 417
rect 703 315 737 349
rect 797 443 831 477
rect 797 375 831 409
rect 797 307 831 341
rect 891 455 925 489
rect 891 357 925 391
rect 985 443 1019 477
rect 985 375 1019 409
rect 985 307 1019 341
rect 1079 455 1113 489
rect 1079 357 1113 391
rect 1173 443 1207 477
rect 1173 375 1207 409
rect 1173 307 1207 341
rect 1267 455 1301 489
rect 1267 357 1301 391
rect 1361 443 1395 477
rect 1361 375 1395 409
rect 1361 307 1395 341
rect 1455 445 1489 479
rect 1455 377 1489 411
rect 1455 309 1489 343
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 749 497 785 523
rect 843 497 879 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1125 497 1161 523
rect 1219 497 1255 523
rect 1313 497 1349 523
rect 1407 497 1443 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 749 282 785 297
rect 843 282 879 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1125 282 1161 297
rect 1219 282 1255 297
rect 1313 282 1349 297
rect 1407 282 1443 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 747 265 787 282
rect 841 265 881 282
rect 935 265 975 282
rect 1029 265 1069 282
rect 1123 265 1163 282
rect 1217 265 1257 282
rect 1311 265 1351 282
rect 1405 265 1445 282
rect 65 249 131 265
rect 65 215 81 249
rect 115 215 131 249
rect 65 199 131 215
rect 173 249 307 265
rect 173 215 189 249
rect 223 215 257 249
rect 291 215 307 249
rect 173 199 307 215
rect 349 249 403 265
rect 349 215 359 249
rect 393 215 403 249
rect 349 199 403 215
rect 455 249 639 265
rect 455 215 589 249
rect 623 215 639 249
rect 455 199 639 215
rect 747 249 1456 265
rect 747 215 769 249
rect 803 215 837 249
rect 871 215 905 249
rect 939 215 973 249
rect 1007 215 1041 249
rect 1075 215 1109 249
rect 1143 215 1177 249
rect 1211 215 1456 249
rect 747 199 1456 215
rect 101 177 131 199
rect 183 177 213 199
rect 267 177 297 199
rect 349 177 379 199
rect 465 177 495 199
rect 549 177 579 199
rect 757 177 787 199
rect 841 177 871 199
rect 945 177 975 199
rect 1029 177 1059 199
rect 1133 177 1163 199
rect 1217 177 1247 199
rect 1321 177 1351 199
rect 1405 177 1435 199
rect 101 21 131 47
rect 183 21 213 47
rect 267 21 297 47
rect 349 21 379 47
rect 465 21 495 47
rect 549 21 579 47
rect 757 21 787 47
rect 841 21 871 47
rect 945 21 975 47
rect 1029 21 1059 47
rect 1133 21 1163 47
rect 1217 21 1247 47
rect 1321 21 1351 47
rect 1405 21 1435 47
<< polycont >>
rect 81 215 115 249
rect 189 215 223 249
rect 257 215 291 249
rect 359 215 393 249
rect 589 215 623 249
rect 769 215 803 249
rect 837 215 871 249
rect 905 215 939 249
rect 973 215 1007 249
rect 1041 215 1075 249
rect 1109 215 1143 249
rect 1177 215 1211 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 19 485 85 493
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 119 478 173 527
rect 119 444 129 478
rect 163 444 173 478
rect 119 428 173 444
rect 207 477 273 493
rect 207 443 223 477
rect 257 443 273 477
rect 19 383 35 417
rect 69 394 85 417
rect 207 394 273 443
rect 307 478 361 527
rect 307 444 317 478
rect 351 444 361 478
rect 307 428 361 444
rect 395 485 649 493
rect 395 479 599 485
rect 395 445 411 479
rect 445 459 599 479
rect 445 445 455 459
rect 395 411 455 445
rect 583 451 599 459
rect 633 451 649 485
rect 395 394 411 411
rect 69 383 223 394
rect 19 360 223 383
rect 257 377 411 394
rect 445 377 455 411
rect 257 360 455 377
rect 19 349 71 360
rect 19 315 35 349
rect 69 315 71 349
rect 409 343 455 360
rect 19 292 71 315
rect 105 292 375 326
rect 409 309 411 343
rect 445 309 455 343
rect 409 292 455 309
rect 489 409 549 425
rect 489 375 505 409
rect 539 375 549 409
rect 489 358 549 375
rect 583 391 649 451
rect 489 341 539 358
rect 583 357 599 391
rect 633 357 649 391
rect 697 485 747 527
rect 697 451 703 485
rect 737 451 747 485
rect 697 417 747 451
rect 697 383 703 417
rect 737 383 747 417
rect 489 307 505 341
rect 697 349 747 383
rect 105 258 139 292
rect 341 258 375 292
rect 19 249 139 258
rect 19 215 81 249
rect 115 215 139 249
rect 19 211 139 215
rect 173 249 307 258
rect 173 215 189 249
rect 223 215 257 249
rect 291 215 307 249
rect 173 211 307 215
rect 341 249 409 258
rect 341 215 359 249
rect 393 215 409 249
rect 341 211 409 215
rect 489 177 539 307
rect 573 249 639 323
rect 697 315 703 349
rect 737 315 747 349
rect 697 299 747 315
rect 787 477 841 493
rect 787 443 797 477
rect 831 443 841 477
rect 787 409 841 443
rect 787 375 797 409
rect 831 375 841 409
rect 787 341 841 375
rect 875 489 941 527
rect 875 455 891 489
rect 925 455 941 489
rect 875 391 941 455
rect 875 357 891 391
rect 925 357 941 391
rect 975 477 1029 493
rect 975 443 985 477
rect 1019 443 1029 477
rect 975 409 1029 443
rect 975 375 985 409
rect 1019 375 1029 409
rect 787 307 797 341
rect 831 323 841 341
rect 975 341 1029 375
rect 1063 489 1129 527
rect 1063 455 1079 489
rect 1113 455 1129 489
rect 1063 391 1129 455
rect 1063 357 1079 391
rect 1113 357 1129 391
rect 1163 477 1217 493
rect 1163 443 1173 477
rect 1207 443 1217 477
rect 1163 409 1217 443
rect 1163 375 1173 409
rect 1207 375 1217 409
rect 975 323 985 341
rect 831 307 985 323
rect 1019 323 1029 341
rect 1163 341 1217 375
rect 1251 489 1317 527
rect 1251 455 1267 489
rect 1301 455 1317 489
rect 1251 391 1317 455
rect 1251 357 1267 391
rect 1301 357 1317 391
rect 1351 477 1405 493
rect 1351 443 1361 477
rect 1395 443 1405 477
rect 1351 409 1405 443
rect 1351 375 1361 409
rect 1395 375 1405 409
rect 1163 323 1173 341
rect 1019 307 1173 323
rect 1207 323 1217 341
rect 1351 341 1405 375
rect 1351 323 1361 341
rect 1207 307 1361 323
rect 1395 307 1405 341
rect 787 289 1405 307
rect 1443 479 1505 527
rect 1443 445 1455 479
rect 1489 445 1505 479
rect 1443 411 1505 445
rect 1443 377 1455 411
rect 1489 377 1505 411
rect 1443 343 1505 377
rect 1443 309 1455 343
rect 1489 309 1505 343
rect 1443 289 1505 309
rect 573 215 589 249
rect 623 215 639 249
rect 573 211 639 215
rect 713 249 1227 255
rect 713 215 769 249
rect 803 215 837 249
rect 871 215 905 249
rect 939 215 973 249
rect 1007 215 1041 249
rect 1075 215 1109 249
rect 1143 215 1177 249
rect 1211 215 1227 249
rect 713 207 1227 215
rect 713 177 747 207
rect 41 161 107 177
rect 41 127 57 161
rect 91 127 107 161
rect 41 93 107 127
rect 41 59 57 93
rect 91 59 107 93
rect 41 17 107 59
rect 207 169 747 177
rect 1309 173 1359 289
rect 207 165 505 169
rect 207 131 223 165
rect 257 135 505 165
rect 539 135 747 169
rect 781 165 1411 173
rect 257 131 273 135
rect 207 93 273 131
rect 489 101 549 135
rect 781 131 797 165
rect 831 139 985 165
rect 831 131 847 139
rect 207 59 223 93
rect 257 59 273 93
rect 207 55 273 59
rect 389 93 455 101
rect 389 59 405 93
rect 439 59 455 93
rect 389 17 455 59
rect 489 67 505 101
rect 539 67 549 101
rect 489 51 549 67
rect 583 93 747 101
rect 583 59 599 93
rect 633 59 697 93
rect 731 59 747 93
rect 583 17 747 59
rect 781 89 847 131
rect 969 131 985 139
rect 1019 139 1173 165
rect 1019 131 1035 139
rect 781 55 797 89
rect 831 55 847 89
rect 781 51 847 55
rect 881 89 935 105
rect 881 55 891 89
rect 925 55 935 89
rect 881 17 935 55
rect 969 89 1035 131
rect 1157 131 1173 139
rect 1207 139 1361 165
rect 1207 131 1223 139
rect 969 55 985 89
rect 1019 55 1035 89
rect 969 51 1035 55
rect 1069 89 1123 105
rect 1069 55 1079 89
rect 1113 55 1123 89
rect 1069 17 1123 55
rect 1157 89 1223 131
rect 1345 131 1361 139
rect 1395 131 1411 165
rect 1157 55 1173 89
rect 1207 55 1223 89
rect 1157 51 1223 55
rect 1257 89 1311 105
rect 1257 55 1267 89
rect 1301 55 1311 89
rect 1257 17 1311 55
rect 1345 89 1411 131
rect 1345 55 1361 89
rect 1395 55 1411 89
rect 1345 51 1411 55
rect 1445 165 1495 181
rect 1479 131 1495 165
rect 1445 89 1495 131
rect 1479 55 1495 89
rect 1445 17 1495 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a21o_8
flabel locali s 29 221 63 255 0 FreeSans 200 180 0 0 A2
port 2 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 200 180 0 0 A1
port 1 nsew signal input
flabel locali s 1317 221 1351 255 0 FreeSans 200 180 0 0 X
port 8 nsew signal output
flabel locali s 581 221 615 255 0 FreeSans 200 180 0 0 B1
port 3 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 12538
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 134
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
