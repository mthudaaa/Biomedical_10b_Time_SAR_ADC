magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 3718 582
<< pwell >>
rect 79 21 3673 203
rect 29 -17 63 17
<< scnmos >>
rect 167 47 197 177
rect 271 47 301 177
rect 375 47 405 177
rect 489 47 519 177
rect 641 47 671 177
rect 735 47 765 177
rect 829 47 859 177
rect 923 47 953 177
rect 1017 47 1047 177
rect 1111 47 1141 177
rect 1205 47 1235 177
rect 1299 47 1329 177
rect 1393 47 1423 177
rect 1487 47 1517 177
rect 1581 47 1611 177
rect 1675 47 1705 177
rect 1769 47 1799 177
rect 1863 47 1893 177
rect 1957 47 1987 177
rect 2061 47 2091 177
rect 2145 47 2175 177
rect 2239 47 2269 177
rect 2333 47 2363 177
rect 2427 47 2457 177
rect 2521 47 2551 177
rect 2615 47 2645 177
rect 2709 47 2739 177
rect 2803 47 2833 177
rect 2897 47 2927 177
rect 2991 47 3021 177
rect 3085 47 3115 177
rect 3179 47 3209 177
rect 3273 47 3303 177
rect 3367 47 3397 177
rect 3461 47 3491 177
rect 3565 47 3595 177
<< scpmoshvt >>
rect 115 297 151 497
rect 219 297 255 497
rect 323 297 359 497
rect 427 297 463 497
rect 643 297 679 497
rect 737 297 773 497
rect 831 297 867 497
rect 925 297 961 497
rect 1019 297 1055 497
rect 1113 297 1149 497
rect 1207 297 1243 497
rect 1301 297 1337 497
rect 1395 297 1431 497
rect 1489 297 1525 497
rect 1583 297 1619 497
rect 1677 297 1713 497
rect 1771 297 1807 497
rect 1865 297 1901 497
rect 1959 297 1995 497
rect 2053 297 2089 497
rect 2147 297 2183 497
rect 2241 297 2277 497
rect 2335 297 2371 497
rect 2429 297 2465 497
rect 2523 297 2559 497
rect 2617 297 2653 497
rect 2711 297 2747 497
rect 2805 297 2841 497
rect 2899 297 2935 497
rect 2993 297 3029 497
rect 3087 297 3123 497
rect 3181 297 3217 497
rect 3275 297 3311 497
rect 3369 297 3405 497
rect 3463 297 3499 497
rect 3557 297 3593 497
<< ndiff >>
rect 105 163 167 177
rect 105 129 113 163
rect 147 129 167 163
rect 105 95 167 129
rect 105 61 113 95
rect 147 61 167 95
rect 105 47 167 61
rect 197 169 271 177
rect 197 135 217 169
rect 251 135 271 169
rect 197 101 271 135
rect 197 67 217 101
rect 251 67 271 101
rect 197 47 271 67
rect 301 163 375 177
rect 301 129 321 163
rect 355 129 375 163
rect 301 95 375 129
rect 301 61 321 95
rect 355 61 375 95
rect 301 47 375 61
rect 405 169 489 177
rect 405 135 425 169
rect 459 135 489 169
rect 405 101 489 135
rect 405 67 425 101
rect 459 67 489 101
rect 405 47 489 67
rect 519 163 641 177
rect 519 61 529 163
rect 631 61 641 163
rect 519 47 641 61
rect 671 163 735 177
rect 671 129 691 163
rect 725 129 735 163
rect 671 95 735 129
rect 671 61 691 95
rect 725 61 735 95
rect 671 47 735 61
rect 765 95 829 177
rect 765 61 785 95
rect 819 61 829 95
rect 765 47 829 61
rect 859 163 923 177
rect 859 129 879 163
rect 913 129 923 163
rect 859 95 923 129
rect 859 61 879 95
rect 913 61 923 95
rect 859 47 923 61
rect 953 95 1017 177
rect 953 61 973 95
rect 1007 61 1017 95
rect 953 47 1017 61
rect 1047 163 1111 177
rect 1047 129 1067 163
rect 1101 129 1111 163
rect 1047 95 1111 129
rect 1047 61 1067 95
rect 1101 61 1111 95
rect 1047 47 1111 61
rect 1141 95 1205 177
rect 1141 61 1161 95
rect 1195 61 1205 95
rect 1141 47 1205 61
rect 1235 163 1299 177
rect 1235 129 1255 163
rect 1289 129 1299 163
rect 1235 95 1299 129
rect 1235 61 1255 95
rect 1289 61 1299 95
rect 1235 47 1299 61
rect 1329 95 1393 177
rect 1329 61 1349 95
rect 1383 61 1393 95
rect 1329 47 1393 61
rect 1423 163 1487 177
rect 1423 129 1443 163
rect 1477 129 1487 163
rect 1423 95 1487 129
rect 1423 61 1443 95
rect 1477 61 1487 95
rect 1423 47 1487 61
rect 1517 95 1581 177
rect 1517 61 1537 95
rect 1571 61 1581 95
rect 1517 47 1581 61
rect 1611 163 1675 177
rect 1611 129 1631 163
rect 1665 129 1675 163
rect 1611 95 1675 129
rect 1611 61 1631 95
rect 1665 61 1675 95
rect 1611 47 1675 61
rect 1705 95 1769 177
rect 1705 61 1725 95
rect 1759 61 1769 95
rect 1705 47 1769 61
rect 1799 163 1863 177
rect 1799 129 1819 163
rect 1853 129 1863 163
rect 1799 95 1863 129
rect 1799 61 1819 95
rect 1853 61 1863 95
rect 1799 47 1863 61
rect 1893 95 1957 177
rect 1893 61 1913 95
rect 1947 61 1957 95
rect 1893 47 1957 61
rect 1987 163 2061 177
rect 1987 129 2007 163
rect 2041 129 2061 163
rect 1987 95 2061 129
rect 1987 61 2007 95
rect 2041 61 2061 95
rect 1987 47 2061 61
rect 2091 95 2145 177
rect 2091 61 2101 95
rect 2135 61 2145 95
rect 2091 47 2145 61
rect 2175 163 2239 177
rect 2175 129 2195 163
rect 2229 129 2239 163
rect 2175 95 2239 129
rect 2175 61 2195 95
rect 2229 61 2239 95
rect 2175 47 2239 61
rect 2269 95 2333 177
rect 2269 61 2289 95
rect 2323 61 2333 95
rect 2269 47 2333 61
rect 2363 163 2427 177
rect 2363 129 2383 163
rect 2417 129 2427 163
rect 2363 95 2427 129
rect 2363 61 2383 95
rect 2417 61 2427 95
rect 2363 47 2427 61
rect 2457 95 2521 177
rect 2457 61 2477 95
rect 2511 61 2521 95
rect 2457 47 2521 61
rect 2551 163 2615 177
rect 2551 129 2571 163
rect 2605 129 2615 163
rect 2551 95 2615 129
rect 2551 61 2571 95
rect 2605 61 2615 95
rect 2551 47 2615 61
rect 2645 95 2709 177
rect 2645 61 2665 95
rect 2699 61 2709 95
rect 2645 47 2709 61
rect 2739 163 2803 177
rect 2739 129 2759 163
rect 2793 129 2803 163
rect 2739 95 2803 129
rect 2739 61 2759 95
rect 2793 61 2803 95
rect 2739 47 2803 61
rect 2833 95 2897 177
rect 2833 61 2853 95
rect 2887 61 2897 95
rect 2833 47 2897 61
rect 2927 163 2991 177
rect 2927 129 2947 163
rect 2981 129 2991 163
rect 2927 95 2991 129
rect 2927 61 2947 95
rect 2981 61 2991 95
rect 2927 47 2991 61
rect 3021 95 3085 177
rect 3021 61 3041 95
rect 3075 61 3085 95
rect 3021 47 3085 61
rect 3115 163 3179 177
rect 3115 129 3135 163
rect 3169 129 3179 163
rect 3115 95 3179 129
rect 3115 61 3135 95
rect 3169 61 3179 95
rect 3115 47 3179 61
rect 3209 95 3273 177
rect 3209 61 3229 95
rect 3263 61 3273 95
rect 3209 47 3273 61
rect 3303 163 3367 177
rect 3303 129 3323 163
rect 3357 129 3367 163
rect 3303 95 3367 129
rect 3303 61 3323 95
rect 3357 61 3367 95
rect 3303 47 3367 61
rect 3397 95 3461 177
rect 3397 61 3417 95
rect 3451 61 3461 95
rect 3397 47 3461 61
rect 3491 163 3565 177
rect 3491 129 3511 163
rect 3545 129 3565 163
rect 3491 95 3565 129
rect 3491 61 3511 95
rect 3545 61 3565 95
rect 3491 47 3565 61
rect 3595 95 3647 177
rect 3595 61 3605 95
rect 3639 61 3647 95
rect 3595 47 3647 61
<< pdiff >>
rect 61 485 115 497
rect 61 451 69 485
rect 103 451 115 485
rect 61 417 115 451
rect 61 383 69 417
rect 103 383 115 417
rect 61 349 115 383
rect 61 315 69 349
rect 103 315 115 349
rect 61 297 115 315
rect 151 477 219 497
rect 151 443 163 477
rect 197 443 219 477
rect 151 409 219 443
rect 151 375 163 409
rect 197 375 219 409
rect 151 341 219 375
rect 151 307 163 341
rect 197 307 219 341
rect 151 297 219 307
rect 255 485 323 497
rect 255 451 267 485
rect 301 451 323 485
rect 255 415 323 451
rect 255 381 267 415
rect 301 381 323 415
rect 255 345 323 381
rect 255 311 267 345
rect 301 311 323 345
rect 255 297 323 311
rect 359 477 427 497
rect 359 443 371 477
rect 405 443 427 477
rect 359 409 427 443
rect 359 375 371 409
rect 405 375 427 409
rect 359 341 427 375
rect 359 307 371 341
rect 405 307 427 341
rect 359 297 427 307
rect 463 485 531 497
rect 463 451 475 485
rect 509 451 531 485
rect 463 415 531 451
rect 463 381 475 415
rect 509 381 531 415
rect 463 345 531 381
rect 463 311 475 345
rect 509 311 531 345
rect 463 297 531 311
rect 585 477 643 497
rect 585 443 597 477
rect 631 443 643 477
rect 585 409 643 443
rect 585 375 597 409
rect 631 375 643 409
rect 585 341 643 375
rect 585 307 597 341
rect 631 307 643 341
rect 585 297 643 307
rect 679 485 737 497
rect 679 451 691 485
rect 725 451 737 485
rect 679 417 737 451
rect 679 383 691 417
rect 725 383 737 417
rect 679 297 737 383
rect 773 477 831 497
rect 773 443 785 477
rect 819 443 831 477
rect 773 409 831 443
rect 773 375 785 409
rect 819 375 831 409
rect 773 341 831 375
rect 773 307 785 341
rect 819 307 831 341
rect 773 297 831 307
rect 867 485 925 497
rect 867 451 879 485
rect 913 451 925 485
rect 867 417 925 451
rect 867 383 879 417
rect 913 383 925 417
rect 867 297 925 383
rect 961 477 1019 497
rect 961 443 973 477
rect 1007 443 1019 477
rect 961 409 1019 443
rect 961 375 973 409
rect 1007 375 1019 409
rect 961 341 1019 375
rect 961 307 973 341
rect 1007 307 1019 341
rect 961 297 1019 307
rect 1055 485 1113 497
rect 1055 451 1067 485
rect 1101 451 1113 485
rect 1055 417 1113 451
rect 1055 383 1067 417
rect 1101 383 1113 417
rect 1055 297 1113 383
rect 1149 477 1207 497
rect 1149 443 1161 477
rect 1195 443 1207 477
rect 1149 409 1207 443
rect 1149 375 1161 409
rect 1195 375 1207 409
rect 1149 341 1207 375
rect 1149 307 1161 341
rect 1195 307 1207 341
rect 1149 297 1207 307
rect 1243 485 1301 497
rect 1243 451 1255 485
rect 1289 451 1301 485
rect 1243 417 1301 451
rect 1243 383 1255 417
rect 1289 383 1301 417
rect 1243 297 1301 383
rect 1337 477 1395 497
rect 1337 443 1349 477
rect 1383 443 1395 477
rect 1337 409 1395 443
rect 1337 375 1349 409
rect 1383 375 1395 409
rect 1337 341 1395 375
rect 1337 307 1349 341
rect 1383 307 1395 341
rect 1337 297 1395 307
rect 1431 485 1489 497
rect 1431 451 1443 485
rect 1477 451 1489 485
rect 1431 417 1489 451
rect 1431 383 1443 417
rect 1477 383 1489 417
rect 1431 297 1489 383
rect 1525 477 1583 497
rect 1525 443 1537 477
rect 1571 443 1583 477
rect 1525 409 1583 443
rect 1525 375 1537 409
rect 1571 375 1583 409
rect 1525 341 1583 375
rect 1525 307 1537 341
rect 1571 307 1583 341
rect 1525 297 1583 307
rect 1619 485 1677 497
rect 1619 451 1631 485
rect 1665 451 1677 485
rect 1619 417 1677 451
rect 1619 383 1631 417
rect 1665 383 1677 417
rect 1619 297 1677 383
rect 1713 477 1771 497
rect 1713 443 1725 477
rect 1759 443 1771 477
rect 1713 409 1771 443
rect 1713 375 1725 409
rect 1759 375 1771 409
rect 1713 341 1771 375
rect 1713 307 1725 341
rect 1759 307 1771 341
rect 1713 297 1771 307
rect 1807 485 1865 497
rect 1807 451 1819 485
rect 1853 451 1865 485
rect 1807 417 1865 451
rect 1807 383 1819 417
rect 1853 383 1865 417
rect 1807 297 1865 383
rect 1901 477 1959 497
rect 1901 443 1913 477
rect 1947 443 1959 477
rect 1901 409 1959 443
rect 1901 375 1913 409
rect 1947 375 1959 409
rect 1901 341 1959 375
rect 1901 307 1913 341
rect 1947 307 1959 341
rect 1901 297 1959 307
rect 1995 485 2053 497
rect 1995 451 2007 485
rect 2041 451 2053 485
rect 1995 417 2053 451
rect 1995 383 2007 417
rect 2041 383 2053 417
rect 1995 297 2053 383
rect 2089 477 2147 497
rect 2089 443 2101 477
rect 2135 443 2147 477
rect 2089 409 2147 443
rect 2089 375 2101 409
rect 2135 375 2147 409
rect 2089 341 2147 375
rect 2089 307 2101 341
rect 2135 307 2147 341
rect 2089 297 2147 307
rect 2183 409 2241 497
rect 2183 375 2195 409
rect 2229 375 2241 409
rect 2183 341 2241 375
rect 2183 307 2195 341
rect 2229 307 2241 341
rect 2183 297 2241 307
rect 2277 477 2335 497
rect 2277 443 2289 477
rect 2323 443 2335 477
rect 2277 409 2335 443
rect 2277 375 2289 409
rect 2323 375 2335 409
rect 2277 297 2335 375
rect 2371 409 2429 497
rect 2371 375 2383 409
rect 2417 375 2429 409
rect 2371 341 2429 375
rect 2371 307 2383 341
rect 2417 307 2429 341
rect 2371 297 2429 307
rect 2465 477 2523 497
rect 2465 443 2477 477
rect 2511 443 2523 477
rect 2465 409 2523 443
rect 2465 375 2477 409
rect 2511 375 2523 409
rect 2465 297 2523 375
rect 2559 409 2617 497
rect 2559 375 2571 409
rect 2605 375 2617 409
rect 2559 341 2617 375
rect 2559 307 2571 341
rect 2605 307 2617 341
rect 2559 297 2617 307
rect 2653 477 2711 497
rect 2653 443 2665 477
rect 2699 443 2711 477
rect 2653 409 2711 443
rect 2653 375 2665 409
rect 2699 375 2711 409
rect 2653 297 2711 375
rect 2747 409 2805 497
rect 2747 375 2759 409
rect 2793 375 2805 409
rect 2747 341 2805 375
rect 2747 307 2759 341
rect 2793 307 2805 341
rect 2747 297 2805 307
rect 2841 477 2899 497
rect 2841 443 2853 477
rect 2887 443 2899 477
rect 2841 409 2899 443
rect 2841 375 2853 409
rect 2887 375 2899 409
rect 2841 297 2899 375
rect 2935 409 2993 497
rect 2935 375 2947 409
rect 2981 375 2993 409
rect 2935 341 2993 375
rect 2935 307 2947 341
rect 2981 307 2993 341
rect 2935 297 2993 307
rect 3029 477 3087 497
rect 3029 443 3041 477
rect 3075 443 3087 477
rect 3029 409 3087 443
rect 3029 375 3041 409
rect 3075 375 3087 409
rect 3029 297 3087 375
rect 3123 409 3181 497
rect 3123 375 3135 409
rect 3169 375 3181 409
rect 3123 341 3181 375
rect 3123 307 3135 341
rect 3169 307 3181 341
rect 3123 297 3181 307
rect 3217 477 3275 497
rect 3217 443 3229 477
rect 3263 443 3275 477
rect 3217 409 3275 443
rect 3217 375 3229 409
rect 3263 375 3275 409
rect 3217 297 3275 375
rect 3311 409 3369 497
rect 3311 375 3323 409
rect 3357 375 3369 409
rect 3311 341 3369 375
rect 3311 307 3323 341
rect 3357 307 3369 341
rect 3311 297 3369 307
rect 3405 477 3463 497
rect 3405 443 3417 477
rect 3451 443 3463 477
rect 3405 409 3463 443
rect 3405 375 3417 409
rect 3451 375 3463 409
rect 3405 297 3463 375
rect 3499 409 3557 497
rect 3499 375 3511 409
rect 3545 375 3557 409
rect 3499 341 3557 375
rect 3499 307 3511 341
rect 3545 307 3557 341
rect 3499 297 3557 307
rect 3593 477 3649 497
rect 3593 443 3605 477
rect 3639 443 3649 477
rect 3593 409 3649 443
rect 3593 375 3605 409
rect 3639 375 3649 409
rect 3593 297 3649 375
<< ndiffc >>
rect 113 129 147 163
rect 113 61 147 95
rect 217 135 251 169
rect 217 67 251 101
rect 321 129 355 163
rect 321 61 355 95
rect 425 135 459 169
rect 425 67 459 101
rect 529 61 631 163
rect 691 129 725 163
rect 691 61 725 95
rect 785 61 819 95
rect 879 129 913 163
rect 879 61 913 95
rect 973 61 1007 95
rect 1067 129 1101 163
rect 1067 61 1101 95
rect 1161 61 1195 95
rect 1255 129 1289 163
rect 1255 61 1289 95
rect 1349 61 1383 95
rect 1443 129 1477 163
rect 1443 61 1477 95
rect 1537 61 1571 95
rect 1631 129 1665 163
rect 1631 61 1665 95
rect 1725 61 1759 95
rect 1819 129 1853 163
rect 1819 61 1853 95
rect 1913 61 1947 95
rect 2007 129 2041 163
rect 2007 61 2041 95
rect 2101 61 2135 95
rect 2195 129 2229 163
rect 2195 61 2229 95
rect 2289 61 2323 95
rect 2383 129 2417 163
rect 2383 61 2417 95
rect 2477 61 2511 95
rect 2571 129 2605 163
rect 2571 61 2605 95
rect 2665 61 2699 95
rect 2759 129 2793 163
rect 2759 61 2793 95
rect 2853 61 2887 95
rect 2947 129 2981 163
rect 2947 61 2981 95
rect 3041 61 3075 95
rect 3135 129 3169 163
rect 3135 61 3169 95
rect 3229 61 3263 95
rect 3323 129 3357 163
rect 3323 61 3357 95
rect 3417 61 3451 95
rect 3511 129 3545 163
rect 3511 61 3545 95
rect 3605 61 3639 95
<< pdiffc >>
rect 69 451 103 485
rect 69 383 103 417
rect 69 315 103 349
rect 163 443 197 477
rect 163 375 197 409
rect 163 307 197 341
rect 267 451 301 485
rect 267 381 301 415
rect 267 311 301 345
rect 371 443 405 477
rect 371 375 405 409
rect 371 307 405 341
rect 475 451 509 485
rect 475 381 509 415
rect 475 311 509 345
rect 597 443 631 477
rect 597 375 631 409
rect 597 307 631 341
rect 691 451 725 485
rect 691 383 725 417
rect 785 443 819 477
rect 785 375 819 409
rect 785 307 819 341
rect 879 451 913 485
rect 879 383 913 417
rect 973 443 1007 477
rect 973 375 1007 409
rect 973 307 1007 341
rect 1067 451 1101 485
rect 1067 383 1101 417
rect 1161 443 1195 477
rect 1161 375 1195 409
rect 1161 307 1195 341
rect 1255 451 1289 485
rect 1255 383 1289 417
rect 1349 443 1383 477
rect 1349 375 1383 409
rect 1349 307 1383 341
rect 1443 451 1477 485
rect 1443 383 1477 417
rect 1537 443 1571 477
rect 1537 375 1571 409
rect 1537 307 1571 341
rect 1631 451 1665 485
rect 1631 383 1665 417
rect 1725 443 1759 477
rect 1725 375 1759 409
rect 1725 307 1759 341
rect 1819 451 1853 485
rect 1819 383 1853 417
rect 1913 443 1947 477
rect 1913 375 1947 409
rect 1913 307 1947 341
rect 2007 451 2041 485
rect 2007 383 2041 417
rect 2101 443 2135 477
rect 2101 375 2135 409
rect 2101 307 2135 341
rect 2195 375 2229 409
rect 2195 307 2229 341
rect 2289 443 2323 477
rect 2289 375 2323 409
rect 2383 375 2417 409
rect 2383 307 2417 341
rect 2477 443 2511 477
rect 2477 375 2511 409
rect 2571 375 2605 409
rect 2571 307 2605 341
rect 2665 443 2699 477
rect 2665 375 2699 409
rect 2759 375 2793 409
rect 2759 307 2793 341
rect 2853 443 2887 477
rect 2853 375 2887 409
rect 2947 375 2981 409
rect 2947 307 2981 341
rect 3041 443 3075 477
rect 3041 375 3075 409
rect 3135 375 3169 409
rect 3135 307 3169 341
rect 3229 443 3263 477
rect 3229 375 3263 409
rect 3323 375 3357 409
rect 3323 307 3357 341
rect 3417 443 3451 477
rect 3417 375 3451 409
rect 3511 375 3545 409
rect 3511 307 3545 341
rect 3605 443 3639 477
rect 3605 375 3639 409
<< poly >>
rect 115 497 151 523
rect 219 497 255 523
rect 323 497 359 523
rect 427 497 463 523
rect 643 497 679 523
rect 737 497 773 523
rect 831 497 867 523
rect 925 497 961 523
rect 1019 497 1055 523
rect 1113 497 1149 523
rect 1207 497 1243 523
rect 1301 497 1337 523
rect 1395 497 1431 523
rect 1489 497 1525 523
rect 1583 497 1619 523
rect 1677 497 1713 523
rect 1771 497 1807 523
rect 1865 497 1901 523
rect 1959 497 1995 523
rect 2053 497 2089 523
rect 2147 497 2183 523
rect 2241 497 2277 523
rect 2335 497 2371 523
rect 2429 497 2465 523
rect 2523 497 2559 523
rect 2617 497 2653 523
rect 2711 497 2747 523
rect 2805 497 2841 523
rect 2899 497 2935 523
rect 2993 497 3029 523
rect 3087 497 3123 523
rect 3181 497 3217 523
rect 3275 497 3311 523
rect 3369 497 3405 523
rect 3463 497 3499 523
rect 3557 497 3593 523
rect 115 282 151 297
rect 219 282 255 297
rect 323 282 359 297
rect 427 282 463 297
rect 643 282 679 297
rect 737 282 773 297
rect 831 282 867 297
rect 925 282 961 297
rect 1019 282 1055 297
rect 1113 282 1149 297
rect 1207 282 1243 297
rect 1301 282 1337 297
rect 1395 282 1431 297
rect 1489 282 1525 297
rect 1583 282 1619 297
rect 1677 282 1713 297
rect 1771 282 1807 297
rect 1865 282 1901 297
rect 1959 282 1995 297
rect 2053 282 2089 297
rect 2147 282 2183 297
rect 2241 282 2277 297
rect 2335 282 2371 297
rect 2429 282 2465 297
rect 2523 282 2559 297
rect 2617 282 2653 297
rect 2711 282 2747 297
rect 2805 282 2841 297
rect 2899 282 2935 297
rect 2993 282 3029 297
rect 3087 282 3123 297
rect 3181 282 3217 297
rect 3275 282 3311 297
rect 3369 282 3405 297
rect 3463 282 3499 297
rect 3557 282 3593 297
rect 113 265 153 282
rect 217 265 257 282
rect 321 265 361 282
rect 425 265 465 282
rect 641 265 681 282
rect 735 265 775 282
rect 829 265 869 282
rect 923 265 963 282
rect 1017 265 1057 282
rect 1111 265 1151 282
rect 1205 265 1245 282
rect 1299 265 1339 282
rect 1393 265 1433 282
rect 1487 265 1527 282
rect 1581 265 1621 282
rect 1675 265 1715 282
rect 1769 265 1809 282
rect 1863 265 1903 282
rect 1957 265 1997 282
rect 2051 265 2091 282
rect 21 249 519 265
rect 21 215 31 249
rect 65 215 99 249
rect 133 215 519 249
rect 21 199 519 215
rect 167 177 197 199
rect 271 177 301 199
rect 375 177 405 199
rect 489 177 519 199
rect 641 249 2091 265
rect 641 215 657 249
rect 691 215 735 249
rect 769 215 813 249
rect 847 215 891 249
rect 925 215 969 249
rect 1003 215 1037 249
rect 1071 215 1115 249
rect 1149 215 1193 249
rect 1227 215 1271 249
rect 1305 215 1349 249
rect 1383 215 1417 249
rect 1451 215 1495 249
rect 1529 215 1573 249
rect 1607 215 1651 249
rect 1685 215 1729 249
rect 1763 215 1797 249
rect 1831 215 1875 249
rect 1909 215 1953 249
rect 1987 215 2031 249
rect 2065 215 2091 249
rect 641 199 2091 215
rect 641 177 671 199
rect 735 177 765 199
rect 829 177 859 199
rect 923 177 953 199
rect 1017 177 1047 199
rect 1111 177 1141 199
rect 1205 177 1235 199
rect 1299 177 1329 199
rect 1393 177 1423 199
rect 1487 177 1517 199
rect 1581 177 1611 199
rect 1675 177 1705 199
rect 1769 177 1799 199
rect 1863 177 1893 199
rect 1957 177 1987 199
rect 2061 177 2091 199
rect 2145 265 2185 282
rect 2239 265 2279 282
rect 2333 265 2373 282
rect 2427 265 2467 282
rect 2521 265 2561 282
rect 2615 265 2655 282
rect 2709 265 2749 282
rect 2803 265 2843 282
rect 2897 265 2937 282
rect 2991 265 3031 282
rect 3085 265 3125 282
rect 3179 265 3219 282
rect 3273 265 3313 282
rect 3367 265 3407 282
rect 3461 265 3501 282
rect 3555 265 3595 282
rect 2145 249 3595 265
rect 2145 215 2161 249
rect 2195 215 2239 249
rect 2273 215 2317 249
rect 2351 215 2395 249
rect 2429 215 2473 249
rect 2507 215 2541 249
rect 2575 215 2619 249
rect 2653 215 2697 249
rect 2731 215 2775 249
rect 2809 215 2853 249
rect 2887 215 2921 249
rect 2955 215 2999 249
rect 3033 215 3077 249
rect 3111 215 3155 249
rect 3189 215 3233 249
rect 3267 215 3301 249
rect 3335 215 3379 249
rect 3413 215 3457 249
rect 3491 215 3595 249
rect 2145 199 3595 215
rect 2145 177 2175 199
rect 2239 177 2269 199
rect 2333 177 2363 199
rect 2427 177 2457 199
rect 2521 177 2551 199
rect 2615 177 2645 199
rect 2709 177 2739 199
rect 2803 177 2833 199
rect 2897 177 2927 199
rect 2991 177 3021 199
rect 3085 177 3115 199
rect 3179 177 3209 199
rect 3273 177 3303 199
rect 3367 177 3397 199
rect 3461 177 3491 199
rect 3565 177 3595 199
rect 167 21 197 47
rect 271 21 301 47
rect 375 21 405 47
rect 489 21 519 47
rect 641 21 671 47
rect 735 21 765 47
rect 829 21 859 47
rect 923 21 953 47
rect 1017 21 1047 47
rect 1111 21 1141 47
rect 1205 21 1235 47
rect 1299 21 1329 47
rect 1393 21 1423 47
rect 1487 21 1517 47
rect 1581 21 1611 47
rect 1675 21 1705 47
rect 1769 21 1799 47
rect 1863 21 1893 47
rect 1957 21 1987 47
rect 2061 21 2091 47
rect 2145 21 2175 47
rect 2239 21 2269 47
rect 2333 21 2363 47
rect 2427 21 2457 47
rect 2521 21 2551 47
rect 2615 21 2645 47
rect 2709 21 2739 47
rect 2803 21 2833 47
rect 2897 21 2927 47
rect 2991 21 3021 47
rect 3085 21 3115 47
rect 3179 21 3209 47
rect 3273 21 3303 47
rect 3367 21 3397 47
rect 3461 21 3491 47
rect 3565 21 3595 47
<< polycont >>
rect 31 215 65 249
rect 99 215 133 249
rect 657 215 691 249
rect 735 215 769 249
rect 813 215 847 249
rect 891 215 925 249
rect 969 215 1003 249
rect 1037 215 1071 249
rect 1115 215 1149 249
rect 1193 215 1227 249
rect 1271 215 1305 249
rect 1349 215 1383 249
rect 1417 215 1451 249
rect 1495 215 1529 249
rect 1573 215 1607 249
rect 1651 215 1685 249
rect 1729 215 1763 249
rect 1797 215 1831 249
rect 1875 215 1909 249
rect 1953 215 1987 249
rect 2031 215 2065 249
rect 2161 215 2195 249
rect 2239 215 2273 249
rect 2317 215 2351 249
rect 2395 215 2429 249
rect 2473 215 2507 249
rect 2541 215 2575 249
rect 2619 215 2653 249
rect 2697 215 2731 249
rect 2775 215 2809 249
rect 2853 215 2887 249
rect 2921 215 2955 249
rect 2999 215 3033 249
rect 3077 215 3111 249
rect 3155 215 3189 249
rect 3233 215 3267 249
rect 3301 215 3335 249
rect 3379 215 3413 249
rect 3457 215 3491 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3680 561
rect 60 485 103 527
rect 60 451 69 485
rect 60 417 103 451
rect 60 383 69 417
rect 60 349 103 383
rect 60 315 69 349
rect 60 299 103 315
rect 137 477 223 493
rect 137 443 163 477
rect 197 443 223 477
rect 137 409 223 443
rect 137 375 163 409
rect 197 375 223 409
rect 137 341 223 375
rect 137 307 163 341
rect 197 307 223 341
rect 137 299 223 307
rect 17 249 133 265
rect 17 215 31 249
rect 65 215 99 249
rect 17 199 133 215
rect 177 257 223 299
rect 267 485 311 527
rect 301 451 311 485
rect 267 415 311 451
rect 301 381 311 415
rect 267 345 311 381
rect 301 311 311 345
rect 267 291 311 311
rect 345 477 431 493
rect 345 443 371 477
rect 405 443 431 477
rect 345 409 431 443
rect 345 375 371 409
rect 405 375 431 409
rect 345 341 431 375
rect 345 307 371 341
rect 405 307 431 341
rect 345 257 431 307
rect 475 485 534 527
rect 509 451 534 485
rect 475 415 534 451
rect 509 381 534 415
rect 475 345 534 381
rect 509 311 534 345
rect 475 291 534 311
rect 575 477 639 493
rect 575 443 597 477
rect 631 443 639 477
rect 575 409 639 443
rect 575 375 597 409
rect 631 375 639 409
rect 575 341 639 375
rect 683 485 733 527
rect 683 451 691 485
rect 725 451 733 485
rect 683 417 733 451
rect 683 383 691 417
rect 725 383 733 417
rect 683 367 733 383
rect 777 477 827 493
rect 777 443 785 477
rect 819 443 827 477
rect 777 409 827 443
rect 777 375 785 409
rect 819 375 827 409
rect 575 307 597 341
rect 631 333 639 341
rect 777 341 827 375
rect 871 485 921 527
rect 871 451 879 485
rect 913 451 921 485
rect 871 417 921 451
rect 871 383 879 417
rect 913 383 921 417
rect 871 367 921 383
rect 965 477 1015 493
rect 965 443 973 477
rect 1007 443 1015 477
rect 965 409 1015 443
rect 965 375 973 409
rect 1007 375 1015 409
rect 777 333 785 341
rect 631 307 785 333
rect 819 333 827 341
rect 965 341 1015 375
rect 1059 485 1109 527
rect 1059 451 1067 485
rect 1101 451 1109 485
rect 1059 417 1109 451
rect 1059 383 1067 417
rect 1101 383 1109 417
rect 1059 367 1109 383
rect 1153 477 1203 493
rect 1153 443 1161 477
rect 1195 443 1203 477
rect 1153 409 1203 443
rect 1153 375 1161 409
rect 1195 375 1203 409
rect 965 333 973 341
rect 819 307 973 333
rect 1007 333 1015 341
rect 1153 341 1203 375
rect 1247 485 1297 527
rect 1247 451 1255 485
rect 1289 451 1297 485
rect 1247 417 1297 451
rect 1247 383 1255 417
rect 1289 383 1297 417
rect 1247 367 1297 383
rect 1341 477 1391 493
rect 1341 443 1349 477
rect 1383 443 1391 477
rect 1341 409 1391 443
rect 1341 375 1349 409
rect 1383 375 1391 409
rect 1153 333 1161 341
rect 1007 307 1161 333
rect 1195 333 1203 341
rect 1341 341 1391 375
rect 1435 485 1485 527
rect 1435 451 1443 485
rect 1477 451 1485 485
rect 1435 417 1485 451
rect 1435 383 1443 417
rect 1477 383 1485 417
rect 1435 367 1485 383
rect 1529 477 1579 493
rect 1529 443 1537 477
rect 1571 443 1579 477
rect 1529 409 1579 443
rect 1529 375 1537 409
rect 1571 375 1579 409
rect 1341 333 1349 341
rect 1195 307 1349 333
rect 1383 333 1391 341
rect 1529 341 1579 375
rect 1623 485 1673 527
rect 1623 451 1631 485
rect 1665 451 1673 485
rect 1623 417 1673 451
rect 1623 383 1631 417
rect 1665 383 1673 417
rect 1623 367 1673 383
rect 1717 477 1767 493
rect 1717 443 1725 477
rect 1759 443 1767 477
rect 1717 409 1767 443
rect 1717 375 1725 409
rect 1759 375 1767 409
rect 1529 333 1537 341
rect 1383 307 1537 333
rect 1571 333 1579 341
rect 1717 341 1767 375
rect 1811 485 1861 527
rect 1811 451 1819 485
rect 1853 451 1861 485
rect 1811 417 1861 451
rect 1811 383 1819 417
rect 1853 383 1861 417
rect 1811 367 1861 383
rect 1905 477 1955 493
rect 1905 443 1913 477
rect 1947 443 1955 477
rect 1905 409 1955 443
rect 1905 375 1913 409
rect 1947 375 1955 409
rect 1717 333 1725 341
rect 1571 307 1725 333
rect 1759 333 1767 341
rect 1905 341 1955 375
rect 1999 485 2049 527
rect 1999 451 2007 485
rect 2041 451 2049 485
rect 1999 417 2049 451
rect 1999 383 2007 417
rect 2041 383 2049 417
rect 1999 367 2049 383
rect 2093 477 3647 493
rect 2093 443 2101 477
rect 2135 459 2289 477
rect 2135 443 2143 459
rect 2093 409 2143 443
rect 2281 443 2289 459
rect 2323 459 2477 477
rect 2323 443 2331 459
rect 2093 375 2101 409
rect 2135 375 2143 409
rect 1905 333 1913 341
rect 1759 307 1913 333
rect 1947 333 1955 341
rect 2093 341 2143 375
rect 2093 333 2101 341
rect 1947 307 2101 333
rect 2135 307 2143 341
rect 575 291 2143 307
rect 2187 409 2237 425
rect 2187 375 2195 409
rect 2229 375 2237 409
rect 2187 341 2237 375
rect 2281 409 2331 443
rect 2469 443 2477 459
rect 2511 459 2665 477
rect 2511 443 2519 459
rect 2281 375 2289 409
rect 2323 375 2331 409
rect 2281 359 2331 375
rect 2375 409 2425 425
rect 2375 375 2383 409
rect 2417 375 2425 409
rect 2187 307 2195 341
rect 2229 325 2237 341
rect 2375 341 2425 375
rect 2469 409 2519 443
rect 2657 443 2665 459
rect 2699 459 2853 477
rect 2699 443 2707 459
rect 2469 375 2477 409
rect 2511 375 2519 409
rect 2469 359 2519 375
rect 2563 409 2613 425
rect 2563 375 2571 409
rect 2605 375 2613 409
rect 2375 325 2383 341
rect 2229 307 2383 325
rect 2417 325 2425 341
rect 2563 341 2613 375
rect 2657 409 2707 443
rect 2845 443 2853 459
rect 2887 459 3041 477
rect 2887 443 2895 459
rect 2657 375 2665 409
rect 2699 375 2707 409
rect 2657 359 2707 375
rect 2751 409 2801 425
rect 2751 375 2759 409
rect 2793 375 2801 409
rect 2563 325 2571 341
rect 2417 307 2571 325
rect 2605 325 2613 341
rect 2751 341 2801 375
rect 2845 409 2895 443
rect 3033 443 3041 459
rect 3075 459 3229 477
rect 3075 443 3083 459
rect 2845 375 2853 409
rect 2887 375 2895 409
rect 2845 359 2895 375
rect 2939 409 2989 425
rect 2939 375 2947 409
rect 2981 375 2989 409
rect 2751 325 2759 341
rect 2605 307 2759 325
rect 2793 325 2801 341
rect 2939 341 2989 375
rect 3033 409 3083 443
rect 3221 443 3229 459
rect 3263 459 3417 477
rect 3263 443 3271 459
rect 3033 375 3041 409
rect 3075 375 3083 409
rect 3033 359 3083 375
rect 3127 409 3177 425
rect 3127 375 3135 409
rect 3169 375 3177 409
rect 2939 325 2947 341
rect 2793 307 2947 325
rect 2981 325 2989 341
rect 3127 341 3177 375
rect 3221 409 3271 443
rect 3409 443 3417 459
rect 3451 459 3605 477
rect 3451 443 3459 459
rect 3221 375 3229 409
rect 3263 375 3271 409
rect 3221 359 3271 375
rect 3315 409 3365 425
rect 3315 375 3323 409
rect 3357 375 3365 409
rect 3127 325 3135 341
rect 2981 307 3135 325
rect 3169 325 3177 341
rect 3315 341 3365 375
rect 3409 409 3459 443
rect 3597 443 3605 459
rect 3639 443 3647 477
rect 3409 375 3417 409
rect 3451 375 3459 409
rect 3409 359 3459 375
rect 3503 409 3553 425
rect 3503 375 3511 409
rect 3545 375 3553 409
rect 3315 325 3323 341
rect 3169 307 3323 325
rect 3357 325 3365 341
rect 3503 341 3553 375
rect 3597 409 3647 443
rect 3597 375 3605 409
rect 3639 375 3647 409
rect 3597 359 3647 375
rect 3503 325 3511 341
rect 3357 307 3511 325
rect 3545 325 3553 341
rect 3545 307 3661 325
rect 2187 291 3661 307
rect 177 249 2096 257
rect 177 215 657 249
rect 691 215 735 249
rect 769 215 813 249
rect 847 215 891 249
rect 925 215 969 249
rect 1003 215 1037 249
rect 1071 215 1115 249
rect 1149 215 1193 249
rect 1227 215 1271 249
rect 1305 215 1349 249
rect 1383 215 1417 249
rect 1451 215 1495 249
rect 1529 215 1573 249
rect 1607 215 1651 249
rect 1685 215 1729 249
rect 1763 215 1797 249
rect 1831 215 1875 249
rect 1909 215 1953 249
rect 1987 215 2031 249
rect 2065 215 2096 249
rect 2130 249 3520 257
rect 2130 215 2161 249
rect 2195 215 2239 249
rect 2273 215 2317 249
rect 2351 215 2395 249
rect 2429 215 2473 249
rect 2507 215 2541 249
rect 2575 215 2619 249
rect 2653 215 2697 249
rect 2731 215 2775 249
rect 2809 215 2853 249
rect 2887 215 2921 249
rect 2955 215 2999 249
rect 3033 215 3077 249
rect 3111 215 3155 249
rect 3189 215 3233 249
rect 3267 215 3301 249
rect 3335 215 3379 249
rect 3413 215 3457 249
rect 3491 215 3520 249
rect 177 213 477 215
rect 17 51 63 199
rect 217 169 269 213
rect 97 163 173 165
rect 97 129 113 163
rect 147 129 173 163
rect 97 95 173 129
rect 97 61 113 95
rect 147 61 173 95
rect 97 17 173 61
rect 251 135 269 169
rect 217 101 269 135
rect 251 67 269 101
rect 217 51 269 67
rect 313 163 373 179
rect 313 129 321 163
rect 355 129 373 163
rect 313 95 373 129
rect 313 61 321 95
rect 355 61 373 95
rect 313 17 373 61
rect 417 169 477 213
rect 3554 181 3661 291
rect 417 135 425 169
rect 459 135 477 169
rect 417 101 477 135
rect 417 67 425 101
rect 459 67 477 101
rect 417 51 477 67
rect 521 163 631 181
rect 521 61 529 163
rect 521 17 631 61
rect 665 163 3661 181
rect 665 129 691 163
rect 725 145 879 163
rect 725 129 741 145
rect 665 95 741 129
rect 853 129 879 145
rect 913 145 1067 163
rect 913 129 929 145
rect 665 61 691 95
rect 725 61 741 95
rect 665 51 741 61
rect 785 95 819 111
rect 785 17 819 61
rect 853 95 929 129
rect 1041 129 1067 145
rect 1101 145 1255 163
rect 1101 129 1117 145
rect 853 61 879 95
rect 913 61 929 95
rect 853 51 929 61
rect 973 95 1007 111
rect 973 17 1007 61
rect 1041 95 1117 129
rect 1229 129 1255 145
rect 1289 145 1443 163
rect 1289 129 1305 145
rect 1041 61 1067 95
rect 1101 61 1117 95
rect 1041 51 1117 61
rect 1161 95 1195 111
rect 1161 17 1195 61
rect 1229 95 1305 129
rect 1417 129 1443 145
rect 1477 145 1631 163
rect 1477 129 1493 145
rect 1229 61 1255 95
rect 1289 61 1305 95
rect 1229 51 1305 61
rect 1349 95 1383 111
rect 1349 17 1383 61
rect 1417 95 1493 129
rect 1605 129 1631 145
rect 1665 145 1819 163
rect 1665 129 1681 145
rect 1417 61 1443 95
rect 1477 61 1493 95
rect 1417 51 1493 61
rect 1537 95 1571 111
rect 1537 17 1571 61
rect 1605 95 1681 129
rect 1793 129 1819 145
rect 1853 145 2007 163
rect 1853 129 1869 145
rect 1605 61 1631 95
rect 1665 61 1681 95
rect 1605 51 1681 61
rect 1725 95 1759 111
rect 1725 17 1759 61
rect 1793 95 1869 129
rect 1981 129 2007 145
rect 2041 145 2195 163
rect 2041 129 2057 145
rect 1793 61 1819 95
rect 1853 61 1869 95
rect 1793 51 1869 61
rect 1913 95 1947 111
rect 1913 17 1947 61
rect 1981 95 2057 129
rect 2169 129 2195 145
rect 2229 145 2383 163
rect 2229 129 2245 145
rect 1981 61 2007 95
rect 2041 61 2057 95
rect 1981 51 2057 61
rect 2101 95 2135 111
rect 2101 17 2135 61
rect 2169 95 2245 129
rect 2357 129 2383 145
rect 2417 145 2571 163
rect 2417 129 2433 145
rect 2169 61 2195 95
rect 2229 61 2245 95
rect 2169 51 2245 61
rect 2289 95 2323 111
rect 2289 17 2323 61
rect 2357 95 2433 129
rect 2545 129 2571 145
rect 2605 145 2759 163
rect 2605 129 2621 145
rect 2357 61 2383 95
rect 2417 61 2433 95
rect 2357 51 2433 61
rect 2477 95 2511 111
rect 2477 17 2511 61
rect 2545 95 2621 129
rect 2733 129 2759 145
rect 2793 145 2947 163
rect 2793 129 2809 145
rect 2545 61 2571 95
rect 2605 61 2621 95
rect 2545 51 2621 61
rect 2665 95 2699 111
rect 2665 17 2699 61
rect 2733 95 2809 129
rect 2921 129 2947 145
rect 2981 145 3135 163
rect 2981 129 2997 145
rect 2733 61 2759 95
rect 2793 61 2809 95
rect 2733 51 2809 61
rect 2853 95 2887 111
rect 2853 17 2887 61
rect 2921 95 2997 129
rect 3109 129 3135 145
rect 3169 145 3323 163
rect 3169 129 3185 145
rect 2921 61 2947 95
rect 2981 61 2997 95
rect 2921 51 2997 61
rect 3041 95 3075 111
rect 3041 17 3075 61
rect 3109 95 3185 129
rect 3297 129 3323 145
rect 3357 145 3511 163
rect 3357 129 3373 145
rect 3109 61 3135 95
rect 3169 61 3185 95
rect 3109 51 3185 61
rect 3229 95 3263 111
rect 3229 17 3263 61
rect 3297 95 3373 129
rect 3485 129 3511 145
rect 3545 145 3661 163
rect 3545 129 3561 145
rect 3297 61 3323 95
rect 3357 61 3373 95
rect 3297 51 3373 61
rect 3417 95 3451 111
rect 3417 17 3451 61
rect 3485 95 3561 129
rect 3485 61 3511 95
rect 3545 61 3561 95
rect 3485 51 3561 61
rect 3605 95 3659 111
rect 3639 61 3659 95
rect 3605 17 3659 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3680 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3433 527 3467 561
rect 3525 527 3559 561
rect 3617 527 3651 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
<< metal1 >>
rect 0 561 3680 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3680 561
rect 0 496 3680 527
rect 0 17 3680 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3680 17
rect 0 -48 3680 -17
<< labels >>
flabel locali s 59 221 93 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 3584 289 3618 323 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel locali s 2130 215 3520 257 0 FreeSans 400 0 0 0 SLEEP
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sky130_fd_sc_hdll__lpflow_isobufsrc_16
<< properties >>
string FIXED_BBOX 0 0 3680 544
string GDS_END 2984266
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 2958944
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
