magic
tech sky130A
magscale 1 2
timestamp 1723858470
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 1 201 853 203
rect 1917 201 2111 203
rect 1 21 2111 201
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 173 47 203 177
rect 267 47 297 177
rect 361 47 391 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 747 47 777 177
rect 842 47 872 175
rect 931 47 961 175
rect 1015 47 1045 175
rect 1285 47 1315 175
rect 1392 47 1422 175
rect 1519 47 1549 175
rect 1623 47 1653 175
rect 1883 47 1913 175
rect 1993 47 2023 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 834 297 870 497
rect 1089 297 1125 497
rect 1183 297 1219 497
rect 1277 297 1313 497
rect 1384 297 1420 497
rect 1697 297 1733 497
rect 1791 297 1827 497
rect 1885 297 1921 497
rect 1995 297 2031 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 101 173 177
rect 109 67 129 101
rect 163 67 173 101
rect 109 47 173 67
rect 203 93 267 177
rect 203 59 223 93
rect 257 59 267 93
rect 203 47 267 59
rect 297 109 361 177
rect 297 75 317 109
rect 351 75 361 109
rect 297 47 361 75
rect 391 93 455 177
rect 391 59 411 93
rect 445 59 455 93
rect 391 47 455 59
rect 485 101 549 177
rect 485 67 505 101
rect 539 67 549 101
rect 485 47 549 67
rect 579 93 643 177
rect 579 59 599 93
rect 633 59 643 93
rect 579 47 643 59
rect 673 109 747 177
rect 673 75 693 109
rect 727 75 747 109
rect 673 47 747 75
rect 777 175 827 177
rect 1943 175 1993 177
rect 777 93 842 175
rect 777 59 787 93
rect 821 59 842 93
rect 777 47 842 59
rect 872 93 931 175
rect 872 59 887 93
rect 921 59 931 93
rect 872 47 931 59
rect 961 161 1015 175
rect 961 127 971 161
rect 1005 127 1015 161
rect 961 47 1015 127
rect 1045 93 1285 175
rect 1045 59 1055 93
rect 1089 59 1285 93
rect 1045 47 1285 59
rect 1315 93 1392 175
rect 1315 59 1348 93
rect 1382 59 1392 93
rect 1315 47 1392 59
rect 1422 93 1519 175
rect 1422 59 1451 93
rect 1485 59 1519 93
rect 1422 47 1519 59
rect 1549 161 1623 175
rect 1549 127 1569 161
rect 1603 127 1623 161
rect 1549 47 1623 127
rect 1653 93 1883 175
rect 1653 59 1663 93
rect 1697 59 1883 93
rect 1653 47 1883 59
rect 1913 93 1993 175
rect 1913 59 1949 93
rect 1983 59 1993 93
rect 1913 47 1993 59
rect 2023 109 2085 177
rect 2023 75 2043 109
rect 2077 75 2085 109
rect 2023 47 2085 75
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 297 81 383
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 297 175 375
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 409 363 443
rect 305 375 317 409
rect 351 375 363 409
rect 305 297 363 375
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 477 551 497
rect 493 443 505 477
rect 539 443 551 477
rect 493 409 551 443
rect 493 375 505 409
rect 539 375 551 409
rect 493 297 551 375
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 417 645 451
rect 587 383 599 417
rect 633 383 645 417
rect 587 297 645 383
rect 681 477 739 497
rect 681 443 693 477
rect 727 443 739 477
rect 681 409 739 443
rect 681 375 693 409
rect 727 375 739 409
rect 681 297 739 375
rect 775 485 834 497
rect 775 451 787 485
rect 821 451 834 485
rect 775 297 834 451
rect 870 485 1089 497
rect 870 451 942 485
rect 976 451 1089 485
rect 870 297 1089 451
rect 1125 401 1183 497
rect 1125 367 1137 401
rect 1171 367 1183 401
rect 1125 297 1183 367
rect 1219 485 1277 497
rect 1219 451 1231 485
rect 1265 451 1277 485
rect 1219 297 1277 451
rect 1313 485 1384 497
rect 1313 451 1335 485
rect 1369 451 1384 485
rect 1313 297 1384 451
rect 1420 485 1697 497
rect 1420 451 1432 485
rect 1466 451 1697 485
rect 1420 297 1697 451
rect 1733 401 1791 497
rect 1733 367 1745 401
rect 1779 367 1791 401
rect 1733 297 1791 367
rect 1827 485 1885 497
rect 1827 451 1839 485
rect 1873 451 1885 485
rect 1827 297 1885 451
rect 1921 485 1995 497
rect 1921 451 1949 485
rect 1983 451 1995 485
rect 1921 297 1995 451
rect 2031 477 2085 497
rect 2031 443 2043 477
rect 2077 443 2085 477
rect 2031 409 2085 443
rect 2031 375 2043 409
rect 2077 375 2085 409
rect 2031 297 2085 375
<< ndiffc >>
rect 35 59 69 93
rect 129 67 163 101
rect 223 59 257 93
rect 317 75 351 109
rect 411 59 445 93
rect 505 67 539 101
rect 599 59 633 93
rect 693 75 727 109
rect 787 59 821 93
rect 887 59 921 93
rect 971 127 1005 161
rect 1055 59 1089 93
rect 1348 59 1382 93
rect 1451 59 1485 93
rect 1569 127 1603 161
rect 1663 59 1697 93
rect 1949 59 1983 93
rect 2043 75 2077 109
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 129 443 163 477
rect 129 375 163 409
rect 223 451 257 485
rect 223 383 257 417
rect 317 443 351 477
rect 317 375 351 409
rect 411 451 445 485
rect 411 383 445 417
rect 505 443 539 477
rect 505 375 539 409
rect 599 451 633 485
rect 599 383 633 417
rect 693 443 727 477
rect 693 375 727 409
rect 787 451 821 485
rect 942 451 976 485
rect 1137 367 1171 401
rect 1231 451 1265 485
rect 1335 451 1369 485
rect 1432 451 1466 485
rect 1745 367 1779 401
rect 1839 451 1873 485
rect 1949 451 1983 485
rect 2043 443 2077 477
rect 2043 375 2077 409
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 834 497 870 523
rect 1089 497 1125 523
rect 1183 497 1219 523
rect 1277 497 1313 523
rect 1384 497 1420 523
rect 1697 497 1733 523
rect 1791 497 1827 523
rect 1885 497 1921 523
rect 1995 497 2031 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 834 282 870 297
rect 1089 282 1125 297
rect 1183 282 1219 297
rect 1277 282 1313 297
rect 1384 282 1420 297
rect 1697 282 1733 297
rect 1791 282 1827 297
rect 1885 282 1921 297
rect 1995 282 2031 297
rect 79 269 119 282
rect 173 269 213 282
rect 267 269 307 282
rect 361 269 401 282
rect 455 269 495 282
rect 549 269 589 282
rect 643 269 683 282
rect 737 269 777 282
rect 79 249 777 269
rect 832 265 872 282
rect 79 215 233 249
rect 267 215 311 249
rect 345 215 379 249
rect 413 215 457 249
rect 491 215 535 249
rect 569 215 613 249
rect 647 215 691 249
rect 725 215 777 249
rect 79 199 777 215
rect 819 249 884 265
rect 819 215 829 249
rect 863 215 884 249
rect 819 199 884 215
rect 931 249 1045 265
rect 931 215 941 249
rect 975 215 1045 249
rect 79 177 109 199
rect 173 177 203 199
rect 267 177 297 199
rect 361 177 391 199
rect 455 177 485 199
rect 549 177 579 199
rect 643 177 673 199
rect 747 177 777 199
rect 842 175 872 199
rect 931 192 1045 215
rect 1087 249 1221 282
rect 1275 265 1315 282
rect 1382 265 1422 282
rect 1087 215 1116 249
rect 1150 215 1221 249
rect 1087 199 1221 215
rect 1263 249 1327 265
rect 1263 215 1273 249
rect 1307 215 1327 249
rect 1263 199 1327 215
rect 1369 249 1446 265
rect 1369 215 1379 249
rect 1413 215 1446 249
rect 1369 199 1446 215
rect 1515 249 1653 265
rect 1515 215 1525 249
rect 1559 215 1653 249
rect 1515 199 1653 215
rect 1695 249 1829 282
rect 1883 265 1923 282
rect 1993 265 2033 282
rect 1695 215 1785 249
rect 1819 215 1829 249
rect 1695 199 1829 215
rect 1873 249 1937 265
rect 1873 215 1883 249
rect 1917 215 1937 249
rect 1873 199 1937 215
rect 1993 249 2067 265
rect 1993 215 2013 249
rect 2047 215 2067 249
rect 1993 199 2067 215
rect 931 175 961 192
rect 1015 175 1045 192
rect 1285 175 1315 199
rect 1392 175 1422 199
rect 1519 192 1653 199
rect 1519 175 1549 192
rect 1623 175 1653 192
rect 1883 175 1913 199
rect 1993 177 2023 199
rect 79 21 109 47
rect 173 21 203 47
rect 267 21 297 47
rect 361 21 391 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 747 21 777 47
rect 842 21 872 47
rect 931 21 961 47
rect 1015 21 1045 47
rect 1285 21 1315 47
rect 1392 21 1422 47
rect 1519 21 1549 47
rect 1623 21 1653 47
rect 1883 21 1913 47
rect 1993 21 2023 47
<< polycont >>
rect 233 215 267 249
rect 311 215 345 249
rect 379 215 413 249
rect 457 215 491 249
rect 535 215 569 249
rect 613 215 647 249
rect 691 215 725 249
rect 829 215 863 249
rect 941 215 975 249
rect 1116 215 1150 249
rect 1273 215 1307 249
rect 1379 215 1413 249
rect 1525 215 1559 249
rect 1785 215 1819 249
rect 1883 215 1917 249
rect 2013 215 2047 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 18 485 85 527
rect 18 451 35 485
rect 69 451 85 485
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 121 477 163 493
rect 121 443 129 477
rect 121 409 163 443
rect 121 375 129 409
rect 197 485 273 527
rect 197 451 223 485
rect 257 451 273 485
rect 197 417 273 451
rect 197 383 223 417
rect 257 383 273 417
rect 317 477 351 493
rect 317 409 351 443
rect 121 349 163 375
rect 385 485 461 527
rect 385 451 411 485
rect 445 451 461 485
rect 385 417 461 451
rect 385 383 411 417
rect 445 383 461 417
rect 505 477 539 493
rect 505 409 539 443
rect 317 349 351 375
rect 573 485 649 527
rect 573 451 599 485
rect 633 451 649 485
rect 573 417 649 451
rect 573 383 599 417
rect 633 383 649 417
rect 693 477 727 493
rect 761 485 837 527
rect 1335 485 1369 527
rect 1933 485 2009 527
rect 761 451 787 485
rect 821 451 837 485
rect 926 451 942 485
rect 976 451 1231 485
rect 1265 451 1281 485
rect 1406 451 1432 485
rect 1466 451 1839 485
rect 1873 451 1889 485
rect 1933 451 1949 485
rect 1983 451 2009 485
rect 2043 477 2077 493
rect 693 409 727 443
rect 1335 435 1369 451
rect 2043 417 2077 443
rect 505 349 539 375
rect 1883 409 2077 417
rect 693 349 727 375
rect 121 315 727 349
rect 761 367 1137 401
rect 1171 367 1745 401
rect 1779 367 1795 401
rect 1883 383 2043 409
rect 121 161 173 315
rect 761 249 795 367
rect 1883 333 1927 383
rect 2043 359 2077 375
rect 217 215 233 249
rect 267 215 311 249
rect 345 215 379 249
rect 413 215 457 249
rect 491 215 535 249
rect 569 215 613 249
rect 647 215 691 249
rect 725 215 795 249
rect 761 161 795 215
rect 829 323 1317 333
rect 829 299 1234 323
rect 829 249 873 299
rect 1268 289 1317 323
rect 941 255 985 265
rect 863 215 873 249
rect 972 249 985 255
rect 829 199 873 215
rect 975 215 985 249
rect 941 199 985 215
rect 1116 249 1160 265
rect 1150 215 1160 249
rect 121 127 727 161
rect 761 127 971 161
rect 1005 153 1034 161
rect 1005 127 1068 153
rect 1116 163 1160 215
rect 1234 249 1317 289
rect 1234 215 1273 249
rect 1307 215 1317 249
rect 1234 199 1317 215
rect 1379 299 1927 333
rect 1379 249 1423 299
rect 1413 215 1423 249
rect 1525 249 1569 265
rect 1379 199 1423 215
rect 1465 215 1525 233
rect 1559 215 1569 249
rect 1465 199 1569 215
rect 1777 255 1834 265
rect 1811 249 1834 255
rect 1777 215 1785 221
rect 1819 215 1834 249
rect 1777 199 1834 215
rect 1883 249 1927 299
rect 1917 215 1927 249
rect 1465 163 1499 199
rect 1116 129 1499 163
rect 121 101 163 127
rect 18 59 35 93
rect 69 59 85 93
rect 18 17 85 59
rect 121 67 129 101
rect 317 109 351 127
rect 121 51 163 67
rect 197 59 223 93
rect 257 59 273 93
rect 505 101 539 127
rect 317 59 351 75
rect 385 59 411 93
rect 445 59 461 93
rect 197 17 273 59
rect 385 17 461 59
rect 693 109 727 127
rect 505 51 539 67
rect 573 59 599 93
rect 633 59 649 93
rect 693 59 727 75
rect 761 59 787 93
rect 821 59 837 93
rect 871 59 887 93
rect 921 59 1055 93
rect 1089 59 1105 93
rect 1151 85 1278 129
rect 1543 127 1569 161
rect 1603 153 1630 161
rect 1664 153 1674 187
rect 1603 127 1674 153
rect 1883 163 1927 215
rect 1995 289 2047 323
rect 1961 249 2047 289
rect 1961 215 2013 249
rect 1961 199 2047 215
rect 1883 129 2077 163
rect 2043 109 2077 129
rect 1332 59 1348 93
rect 1382 59 1398 93
rect 1435 59 1451 93
rect 1485 59 1663 93
rect 1697 59 1713 93
rect 1933 59 1949 93
rect 1983 59 2009 93
rect 2043 59 2077 75
rect 573 17 649 59
rect 761 17 837 59
rect 1332 17 1398 59
rect 1933 17 2009 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 1234 289 1268 323
rect 938 249 972 255
rect 938 221 941 249
rect 941 221 972 249
rect 1034 153 1068 187
rect 1777 249 1811 255
rect 1777 221 1785 249
rect 1785 221 1811 249
rect 1630 153 1664 187
rect 1961 289 1995 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 1222 323 1280 329
rect 1222 289 1234 323
rect 1268 320 1280 323
rect 1949 323 2007 329
rect 1949 320 1961 323
rect 1268 292 1961 320
rect 1268 289 1280 292
rect 1222 283 1280 289
rect 1949 289 1961 292
rect 1995 289 2007 323
rect 1949 283 2007 289
rect 924 255 992 261
rect 924 221 938 255
rect 972 252 992 255
rect 1753 255 1823 261
rect 1753 252 1777 255
rect 972 224 1777 252
rect 972 221 992 224
rect 924 215 992 221
rect 1753 221 1777 224
rect 1811 221 1823 255
rect 1753 215 1823 221
rect 1022 187 1080 193
rect 1022 153 1034 187
rect 1068 184 1080 187
rect 1618 187 1686 193
rect 1618 184 1630 187
rect 1068 156 1630 184
rect 1068 153 1080 156
rect 1022 147 1080 153
rect 1618 153 1630 156
rect 1664 153 1686 187
rect 1618 147 1686 153
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< labels >>
flabel metal1 s 1961 289 1995 323 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel metal1 s 1777 221 1811 255 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel locali s 1225 85 1259 119 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
rlabel comment s 0 0 0 0 4 mux2_8
<< properties >>
string FIXED_BBOX 0 0 2116 544
string GDS_END 1447258
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_START 1433798
string LEFclass CORE
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
